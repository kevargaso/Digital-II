
module mult_32 (input clk, input \B[7] , input rst, output \pp[5] , input \A[0] , output \pp[30] , output \pp[28] , output \pp[31] , output \pp[29] , output \pp[22] , output \pp[27] , output \pp[26] , output \pp[25] , output \pp[24] , output \pp[23] , input \A[3] , input \B[1] , input \B[0] , input \A[1] , input \A[5] , input \B[2] , input \A[7] , input \B[3] , input \B[4] , output done, input \B[5] , input \B[6] , input init, output \pp[9] , input \A[2] , input \A[4] , input \B[8] , input \B[9] , input \B[13] , input \B[12] , input \A[8] , input \A[12] , input \B[14] , input \B[10] , input \B[11] , output \pp[6] , input \B[15] , output \pp[12] , input \A[15] , input \A[9] , input \A[6] , output \pp[0] , output \pp[1] , output \pp[2] , output \pp[3] , output \pp[4] , output \pp[7] , output \pp[8] , output \pp[10] , output \pp[11] , output \pp[13] , output \pp[14] , output \pp[15] , input \A[14] , input \A[13] , input \A[11] , input \A[10] , output \pp[16] , output \pp[17] , output \pp[18] , output \pp[19] , output \pp[20] , output \pp[21] );

wire n2, n3, clk, \B[7] , rst, \A[0] , \pp[30] , \A[3] , \B[1] , \B[0] ;
wire \A[1] , \A[5] , \B[2] , \A[7] , n27, \B[3] , \B[4] , n34, n38, n42;
wire n43, n44, n45, n46, n48, \B[5] , \B[6] , init, n56, n57;
wire n58, n59, n60, n61, n62, n63, n64, \A[2] , n71, n72;
wire n73, \A[4] , \B[8] , \B[9] , \B[13] , \B[12] , \A[8] , \A[12] , \B[14] , \B[10] ;
wire \B[11] , n99, \B[15] , \A[15] , \A[9] , \A[6] , \A[14] , \A[13] , \A[11] , \A[10] ;
wire n135, n136, n137, n138, n139, n140, n141, n142, n144, n145;
wire n146, n147, n148, n149, n150, n151, n160, n161, n162, n163;
wire n164, n165, n166, n167, n175, n176, n177, n178, n179, n180;
wire n181, n182, n183, n184, n185, n186, n187, n188, n189, n190;
wire n191, n192, n193, n194, n195, n196, n197, n198, n199, n200;
wire n201, n202, n203, n204, n205, n206, n207, n208, n209, n210;
wire n211, n212, n213, n214, n215, n216, n217, n218, n219, n220;
wire n221, n222, n223, n224, n225, n226, n227, n228, n229, n230;
wire n231, n232, n233, n234, n235, n236, n237, n238, n239, n240;
wire n241, n242, n243, n244, n245, n246, n247, n248, n249, n250;
wire n251, n252, n253, n254, n255, n256, n257, n258, n259, n260;
wire n261, n262, n263, n264, n265, n266, n267, n268, n269, n270;
wire n271, n272, n273, n274, n275, n276, n277, n278, n279, n280;
wire n281, n282, n283, n284, n285, n286, n287, n288, n289, n290;
wire n291, n292, n293, n294, n295, n296, n297, n298, n299;
reg n1 = 0, \pp[5]  = 0, \pp[28]  = 0, \pp[31]  = 0, \pp[29]  = 0, \pp[22]  = 0, \pp[27]  = 0, \pp[26]  = 0, \pp[25]  = 0, \pp[24]  = 0;
reg \pp[23]  = 0, n22 = 0, n28 = 0, n29 = 0, n30 = 0, n33 = 0, n35 = 0, n36 = 0, n37 = 0, n39 = 0;
reg n40 = 0, done = 0, n47 = 0, n49 = 0, n50 = 0, n53 = 0, n55 = 0, n65 = 0, n66 = 0, n67 = 0;
reg n68 = 0, \pp[9]  = 0, n75 = 0, n76 = 0, n79 = 0, n80 = 0, n81 = 0, n82 = 0, n87 = 0, n88 = 0;
reg n89 = 0, n90 = 0, n91 = 0, n92 = 0, n93 = 0, n95 = 0, n98 = 0, \pp[6]  = 0, n102 = 0, n103 = 0;
reg n104 = 0, n105 = 0, n106 = 0, \pp[12]  = 0, \pp[0]  = 0, \pp[1]  = 0, \pp[2]  = 0, \pp[3]  = 0, \pp[4]  = 0, \pp[7]  = 0;
reg \pp[8]  = 0, \pp[10]  = 0, \pp[11]  = 0, \pp[13]  = 0, \pp[14]  = 0, \pp[15]  = 0, \pp[16]  = 0, \pp[17]  = 0, \pp[18]  = 0, \pp[19]  = 0;
reg \pp[20]  = 0, \pp[21]  = 0, n133 = 0, n134 = 0, n143 = 0, n152 = 0, n153 = 0, n154 = 0, n155 = 0, n156 = 0;
reg n157 = 0, n158 = 0, n159 = 0, n168 = 0, n169 = 0, n170 = 0, n171 = 0, n172 = 0, n173 = 0, n174 = 0;
assign n223 = 0;
assign n255 = 1;

// Debug Symbols
wire \_w_reset_$glb_sr = n1;
wire \_control0.add_SB_LUT4_I3_O_$glb_ce = n2;
wire \_control0.sh_SB_LUT4_I2_O_$glb_ce = n3;
wire \_clk$SB_IO_IN_$glb_clk = clk;
wire \_B[7]$SB_IO_IN = \B[7] ;
wire \_rst$SB_IO_IN = rst;
wire \_pp[5]$SB_IO_OUT = \pp[5] ;
wire \_A[0]$SB_IO_IN = \A[0] ;
wire \_clk$SB_IO_IN = clk;
wire \_control0.add_SB_LUT4_I3_O = n2;
wire \_pp[30]$SB_IO_OUT = \pp[30] ;
wire \_pp[28]$SB_IO_OUT = \pp[28] ;
wire \_pp[31]$SB_IO_OUT = \pp[31] ;
wire \_pp[29]$SB_IO_OUT = \pp[29] ;
wire \_pp[22]$SB_IO_OUT = \pp[22] ;
wire \_pp[27]$SB_IO_OUT = \pp[27] ;
wire \_pp[26]$SB_IO_OUT = \pp[26] ;
wire \_pp[25]$SB_IO_OUT = \pp[25] ;
wire \_pp[24]$SB_IO_OUT = \pp[24] ;
wire \_pp[23]$SB_IO_OUT = \pp[23] ;
wire \_A[3]$SB_IO_IN = \A[3] ;
wire \_B[1]$SB_IO_IN = \B[1] ;
wire \_B[0]$SB_IO_IN = \B[0] ;
wire \_pp[30]$SB_IO_OUT_ = n22;
wire \_A[1]$SB_IO_IN = \A[1] ;
wire \_A[5]$SB_IO_IN = \A[5] ;
wire \_B[2]$SB_IO_IN = \B[2] ;
wire \_A[7]$SB_IO_IN = \A[7] ;
wire \_control0.done_SB_DFFE_Q_D_SB_LUT4_I3_O = n27;
wire \_w_B[4] = n28;
wire \_w_B[5] = n29;
wire \_w_B[6] = n30;
wire \_B[3]$SB_IO_IN = \B[3] ;
wire \_B[4]$SB_IO_IN = \B[4] ;
wire \_w_B[0] = n33;
wire \_control0.lsb_B_SB_LUT4_I0_O[1] = n34;
wire \_w_B[1] = n35;
wire \_w_B[3] = n36;
wire \_w_B[7] = n37;
wire \_control0.lsb_B_SB_LUT4_I0_O[0] = n38;
wire \_w_B[2] = n39;
wire \_w_sh = n40;
wire \_done$SB_IO_OUT = done;
wire \_control0.done_SB_DFFE_Q_D[0] = n42;
wire \_init_SB_LUT4_I1_O[0] = n43;
wire \_control0.sh_SB_LUT4_I2_O = n3;
wire \_init_SB_LUT4_I1_O_SB_LUT4_I1_O[1] = n44;
wire \_init_SB_LUT4_I1_O_SB_LUT4_I1_O[2] = n45;
wire \_rst_SB_LUT4_I2_O = n46;
wire \_control0.state[0] = n47;
wire \_control0.state_SB_DFFSR_Q_R = n48;
wire \_init_SB_LUT4_I1_O[1] = n49;
wire \_init_SB_LUT4_I1_O[2] = n50;
wire \_w_reset = n1;
wire \_B[5]$SB_IO_IN = \B[5] ;
wire \_B[6]$SB_IO_IN = \B[6] ;
wire \_w_B[8] = n53;
wire \_init$SB_IO_IN = init;
wire \_w_add = n55;
wire \_init_SB_LUT4_I1_O_SB_LUT4_I1_O[0] = n56;
wire \_control0.done_SB_DFFE_Q_D_SB_LUT4_I3_1_O[2] = n57;
wire \_rst_SB_LUT4_I3_O[2] = n58;
wire \_rst_SB_LUT4_I2_O_ = n59;
wire \_control0.lsb_B_SB_LUT4_I0_O[3] = n60;
wire \_control0.count_SB_DFFESR_Q_D[1] = n61;
wire \_control0.count_SB_DFFESR_Q_D[2] = n62;
wire \_control0.count_SB_DFFESR_Q_D[3] = n63;
wire \_rst_SB_LUT4_I3_O[2]_ = n64;
wire \_control0.count[1] = n65;
wire \_control0.count[2] = n66;
wire \_control0.count[3] = n67;
wire \_control0.count[0] = n68;
wire \_pp[9]$SB_IO_OUT = \pp[9] ;
wire \_A[2]$SB_IO_IN = \A[2] ;
wire \_control0.lsb_B_SB_LUT4_I0_O[2] = n71;
wire \_control0.count_SB_CARRY_CI_CO[2] = n72;
wire \_control0.count_SB_CARRY_CI_CO[3] = n73;
wire \_A[4]$SB_IO_IN = \A[4] ;
wire \_w_B[13] = n75;
wire \_w_B[14] = n76;
wire \_B[8]$SB_IO_IN = \B[8] ;
wire \_B[9]$SB_IO_IN = \B[9] ;
wire \_w_B[9] = n79;
wire \_w_B[10] = n80;
wire \_w_B[11] = n81;
wire \_w_B[12] = n82;
wire \_B[13]$SB_IO_IN = \B[13] ;
wire \_B[12]$SB_IO_IN = \B[12] ;
wire \_A[8]$SB_IO_IN = \A[8] ;
wire \_A[12]$SB_IO_IN = \A[12] ;
wire \_w_A[2] = n87;
wire \_w_A[4] = n88;
wire \_w_A[5] = n89;
wire \_w_A[3] = n90;
wire \_w_A[7] = n91;
wire \_w_A[6] = n92;
wire \_w_A[1] = n93;
wire \_B[14]$SB_IO_IN = \B[14] ;
wire \_w_B[15] = n95;
wire \_B[10]$SB_IO_IN = \B[10] ;
wire \_B[11]$SB_IO_IN = \B[11] ;
wire \_w_A[0] = n98;
wire \_rsr0.s_B_SB_DFFNESR_Q_R = n99;
wire \_pp[6]$SB_IO_OUT = \pp[6] ;
wire \_B[15]$SB_IO_IN = \B[15] ;
wire \_w_A[12] = n102;
wire \_w_A[11] = n103;
wire \_w_A[8] = n104;
wire \_w_A[10] = n105;
wire \_w_A[9] = n106;
wire \_pp[12]$SB_IO_OUT = \pp[12] ;
wire \_A[15]$SB_IO_IN = \A[15] ;
wire \_A[9]$SB_IO_IN = \A[9] ;
wire \_A[6]$SB_IO_IN = \A[6] ;
wire \_pp[0]$SB_IO_OUT = \pp[0] ;
wire \_pp[1]$SB_IO_OUT = \pp[1] ;
wire \_pp[2]$SB_IO_OUT = \pp[2] ;
wire \_pp[3]$SB_IO_OUT = \pp[3] ;
wire \_pp[4]$SB_IO_OUT = \pp[4] ;
wire \_pp[7]$SB_IO_OUT = \pp[7] ;
wire \_pp[8]$SB_IO_OUT = \pp[8] ;
wire \_pp[10]$SB_IO_OUT = \pp[10] ;
wire \_pp[11]$SB_IO_OUT = \pp[11] ;
wire \_pp[13]$SB_IO_OUT = \pp[13] ;
wire \_pp[14]$SB_IO_OUT = \pp[14] ;
wire \_pp[15]$SB_IO_OUT = \pp[15] ;
wire \_A[14]$SB_IO_IN = \A[14] ;
wire \_A[13]$SB_IO_IN = \A[13] ;
wire \_A[11]$SB_IO_IN = \A[11] ;
wire \_A[10]$SB_IO_IN = \A[10] ;
wire \_pp[16]$SB_IO_OUT = \pp[16] ;
wire \_pp[17]$SB_IO_OUT = \pp[17] ;
wire \_pp[18]$SB_IO_OUT = \pp[18] ;
wire \_pp[19]$SB_IO_OUT = \pp[19] ;
wire \_pp[20]$SB_IO_OUT = \pp[20] ;
wire \_pp[21]$SB_IO_OUT = \pp[21] ;
wire \_w_A[14] = n133;
wire \_w_A[13] = n134;
wire \_acc0.pp_SB_CARRY_I1_CO[1] = n135;
wire \_acc0.pp_SB_CARRY_I1_CO[2] = n136;
wire \_acc0.pp_SB_CARRY_I1_CO[3] = n137;
wire \_acc0.pp_SB_CARRY_I1_CO[4] = n138;
wire \_acc0.pp_SB_CARRY_I1_CO[5] = n139;
wire \_acc0.pp_SB_CARRY_I1_CO[6] = n140;
wire \_acc0.pp_SB_CARRY_I1_CO[7] = n141;
wire \_acc0.pp_SB_CARRY_I1_CO[8] = n142;
wire \_w_A[15] = n143;
wire \_acc0.pp_SB_CARRY_I1_CO[9] = n144;
wire \_acc0.pp_SB_CARRY_I1_CO[10] = n145;
wire \_acc0.pp_SB_CARRY_I1_CO[11] = n146;
wire \_acc0.pp_SB_CARRY_I1_CO[12] = n147;
wire \_acc0.pp_SB_CARRY_I1_CO[13] = n148;
wire \_acc0.pp_SB_CARRY_I1_CO[14] = n149;
wire \_acc0.pp_SB_CARRY_I1_CO[15] = n150;
wire \_acc0.pp_SB_CARRY_I1_CO[16] = n151;
wire \_w_A[21] = n152;
wire \_w_A[20] = n153;
wire \_w_A[18] = n154;
wire \_w_A[19] = n155;
wire \_w_A[16] = n156;
wire \_w_A[22] = n157;
wire \_w_A[23] = n158;
wire \_w_A[17] = n159;
wire \_acc0.pp_SB_CARRY_I1_CO[17] = n160;
wire \_acc0.pp_SB_CARRY_I1_CO[18] = n161;
wire \_acc0.pp_SB_CARRY_I1_CO[19] = n162;
wire \_acc0.pp_SB_CARRY_I1_CO[20] = n163;
wire \_acc0.pp_SB_CARRY_I1_CO[21] = n164;
wire \_acc0.pp_SB_CARRY_I1_CO[22] = n165;
wire \_acc0.pp_SB_CARRY_I1_CO[23] = n166;
wire \_acc0.pp_SB_CARRY_I1_CO[24] = n167;
wire \_w_A[28] = n168;
wire \_w_A[26] = n169;
wire \_w_A[24] = n170;
wire \_w_A[29] = n171;
wire \_w_A[27] = n172;
wire \_w_A[30] = n173;
wire \_w_A[25] = n174;
wire \_acc0.pp_SB_CARRY_I1_CO[25] = n175;
wire \_acc0.pp_SB_CARRY_I1_CO[26] = n176;
wire \_acc0.pp_SB_CARRY_I1_CO[27] = n177;
wire \_acc0.pp_SB_CARRY_I1_CO[28] = n178;
wire \_acc0.pp_SB_CARRY_I1_CO[29] = n179;
wire \_acc0.pp_SB_CARRY_I1_CO[30] = n180;
wire \_acc0.pp_SB_CARRY_I1_CO[31] = n181;

assign n254 = /* LUT    7  2  0 */ 1'b0;
assign n183 = /* LUT   10  3  3 */ (\A[11]  ? (n1 ? 1'b1 : n105) : (n1 ? 1'b0 : n105));
assign n184 = /* LUT    5  2  7 */ (\B[2]  ? (n1 ? 1'b1 : n36) : (n1 ? 1'b0 : n36));
assign n185 = /* LUT    7  2  3 */ (n73 ? !n67 : n67);
assign n186 = /* LUT   11  3  4 */ (n163 ? (n153 ? \pp[20]  : !\pp[20] ) : (n153 ? !\pp[20]  : \pp[20] ));
assign n187 = /* LUT   10  1  6 */ (n89 ? (\A[6]  ? 1'b1 : !n1) : (\A[6]  ? n1 : 1'b0));
assign n188 = /* LUT    5  2  1 */ (n35 ? 1'b0 : (n39 ? 1'b0 : (n33 ? 1'b0 : !n36)));
assign n189 = /* LUT   11  3  6 */ (n165 ? (n157 ? \pp[22]  : !\pp[22] ) : (n157 ? !\pp[22]  : \pp[22] ));
assign n190 = /* LUT    7  2  1 */ (n68 ? !n65 : n65);
assign n191 = /* LUT   10  1  4 */ (n1 ? \A[3]  : n87);
assign n192 = /* LUT   10  1  2 */ (\A[4]  ? (n90 ? 1'b1 : n1) : (n90 ? !n1 : 1'b0));
assign n193 = /* LUT   12  2  4 */ (\A[15]  ? (n1 ? 1'b1 : n133) : (n1 ? 1'b0 : n133));
assign n194 = /* LUT    9  1  1 */ (n1 ? \B[13]  : n76);
assign n195 = /* LUT    1 25  4 */ n22;
assign n196 = /* LUT   12  4  6 */ n171;
assign n197 = /* LUT   10  1  0 */ (n1 ? \A[2]  : n93);
assign n198 = /* LUT    9  1  3 */ (n1 ? \B[14]  : n95);
assign n199 = /* LUT   12  4  4 */ n168;
assign n200 = /* LUT    7  3  4 */ n62;
assign n201 = /* LUT   10  2  6 */ \B[15] ;
assign n202 = /* LUT   12  4  2 */ n174;
assign n203 = /* LUT    7  3  6 */ n63;
assign n204 = /* LUT   10  2  4 */ !n1;
assign n205 = /* LUT    5  3  0 */ (n49 ? (n50 ? 1'b1 : n47) : (n50 ? !n47 : 1'b0));
assign n206 = /* LUT    6  3  1 */ (n49 ? (n50 ? 1'b1 : n47) : (n50 ? 1'b0 : !n47));
assign n207 = /* LUT    5  3  6 */ (n49 ? (n47 ? 1'b0 : !n50) : 1'b0);
assign n208 = /* LUT   11  1  6 */ (n140 ? (\pp[6]  ? n92 : !n92) : (\pp[6]  ? !n92 : n92));
assign n209 = /* LUT    7  3  2 */ n58;
assign n210 = /* LUT    5  3  4 */ n42;
assign n211 = /* LUT   11  1  4 */ (n138 ? (n88 ? \pp[4]  : !\pp[4] ) : (n88 ? !\pp[4]  : \pp[4] ));
assign n212 = /* LUT   11  2  2 */ (n145 ? (\pp[10]  ? n105 : !n105) : (\pp[10]  ? !n105 : n105));
assign n213 = /* LUT    6  3  5 */ (n50 ? (n49 ? 1'b1 : n47) : (n49 ? n47 : 1'b0));
assign n214 = /* LUT   12  1  5 */ (n102 ? (n1 ? \A[13]  : 1'b1) : (n1 ? \A[13]  : 1'b0));
assign n215 = /* LUT    9  2  0 */ (n1 ? \B[9]  : n80);
assign n216 = /* LUT    6  4  4 */ (n49 ? n58 : (n58 ? 1'b1 : !rst));
assign n217 = /* LUT   11  1  2 */ (n136 ? (n87 ? \pp[2]  : !\pp[2] ) : (n87 ? !\pp[2]  : \pp[2] ));
assign n218 = /* LUT   11  2  0 */ (n142 ? (n104 ? \pp[8]  : !\pp[8] ) : (n104 ? !\pp[8]  : \pp[8] ));
assign n219 = /* LUT    6  3  7 */ (n62 ? (n42 ? !n63 : 1'b0) : (n42 ? (n61 ? !n63 : 1'b1) : 1'b0));
assign n220 = /* LUT    5  1  7 */ (n1 ? \B[6]  : n37);
assign n221 = /* LUT    9  2  2 */ (n82 ? 1'b0 : (n95 ? 1'b0 : (n76 ? 1'b0 : !n75)));
assign n222 = /* LUT   11  1  0 */ (\pp[0]  ? !n98 : n98);
assign n224 = /* LUT   11  2  6 */ (n149 ? (n133 ? \pp[14]  : !\pp[14] ) : (n133 ? !\pp[14]  : \pp[14] ));
assign n225 = /* LUT    6  4  0 */ (n50 ? 1'b0 : (n47 ? 1'b0 : !rst));
assign n226 = /* LUT    9  2  4 */ (n81 ? (n1 ? \B[10]  : 1'b1) : (n1 ? \B[10]  : 1'b0));
assign n227 = /* LUT   11  2  4 */ (n147 ? (\pp[12]  ? n102 : !n102) : (\pp[12]  ? !n102 : n102));
assign n228 = /* LUT    5  4  3 */ (n45 ? 1'b1 : (n44 ? !n56 : 1'b0));
assign n229 = /* LUT    6  4  2 */ (n1 ? 1'b1 : n55);
assign n230 = /* LUT    9  2  6 */ (n82 ? (n1 ? \B[11]  : 1'b1) : (n1 ? \B[11]  : 1'b0));
assign n231 = /* LUT    6  2  0 */ (n1 ? 1'b1 : n40);
assign n232 = /* LUT    5  4  1 */ (n49 ? 1'b0 : (n43 ? 1'b0 : !n50));
assign n233 = /* LUT   12  3  6 */ n157;
assign n234 = /* LUT   11  4  5 */ (n179 ? (n171 ? \pp[29]  : !\pp[29] ) : (n171 ? !\pp[29]  : \pp[29] ));
assign n235 = /* LUT   10  3  4 */ (n91 ? (\A[8]  ? 1'b1 : !n1) : (\A[8]  ? n1 : 1'b0));
assign n236 = /* LUT    5  4  7 */ (n49 ? 1'b0 : n47);
assign n237 = /* LUT    9  3  3 */ (n81 ? 1'b0 : (n80 ? 1'b0 : (n53 ? 1'b0 : !n79)));
assign n238 = /* LUT   12  3  4 */ n143;
assign n239 = /* LUT   11  4  7 */ (n181 ? !\pp[31]  : \pp[31] );
assign n240 = /* LUT   10  3  6 */ (n1 ? \A[10]  : n106);
assign n241 = /* LUT   12  3  2 */ n159;
assign n242 = /* LUT   11  3  1 */ (n160 ? (\pp[17]  ? n159 : !n159) : (\pp[17]  ? !n159 : n159));
assign n243 = /* LUT   11  4  1 */ (n175 ? (n174 ? \pp[25]  : !\pp[25] ) : (n174 ? !\pp[25]  : \pp[25] ));
assign n244 = /* LUT    5  2  4 */ (n1 ? \B[3]  : n28);
assign n245 = /* LUT   12  3  0 */ n153;
assign n246 = /* LUT   11  3  3 */ (n162 ? (n155 ? \pp[19]  : !\pp[19] ) : (n155 ? !\pp[19]  : \pp[19] ));
assign n247 = /* LUT   11  4  3 */ (n177 ? (n172 ? \pp[27]  : !\pp[27] ) : (n172 ? !\pp[27]  : \pp[27] ));
assign n248 = /* LUT    5  2  6 */ (n37 ? 1'b0 : (n29 ? 1'b0 : (n28 ? 1'b0 : !n30)));
assign n249 = /* LUT    7  2  2 */ (n72 ? !n66 : n66);
assign n250 = /* LUT   11  3  5 */ (n164 ? (\pp[21]  ? n152 : !n152) : (\pp[21]  ? !n152 : n152));
assign n251 = /* LUT    5  2  0 */ (\B[0]  ? (n35 ? 1'b1 : n1) : (n35 ? !n1 : 1'b0));
assign n252 = /* LUT   11  3  7 */ (n166 ? (\pp[23]  ? n158 : !n158) : (\pp[23]  ? !n158 : n158));
assign n256 = /* LUT   10  1  7 */ (n98 ? (\A[1]  ? 1'b1 : !n1) : (\A[1]  ? n1 : 1'b0));
assign n257 = /* LUT    5  2  2 */ (n1 ? \B[1]  : n39);
assign n258 = /* LUT   10  1  5 */ (\A[7]  ? (n92 ? 1'b1 : n1) : (n92 ? !n1 : 1'b0));
assign n259 = /* LUT   12  4  7 */ n170;
assign n260 = /* LUT   10  1  3 */ (n88 ? (n1 ? \A[5]  : 1'b1) : (n1 ? \A[5]  : 1'b0));
assign n261 = /* LUT   10  2  1 */ \A[0] ;
assign n262 = /* LUT   12  4  5 */ n169;
assign n263 = /* LUT   12  4  3 */ n158;
assign n264 = /* LUT    7  3  7 */ !n68;
assign n265 = /* LUT   12  4  1 */ n172;
assign n266 = /* LUT    5  3  7 */ (init ? (n33 ? 1'b0 : n47) : (n33 ? !n47 : 1'b1));
assign n267 = /* LUT   11  1  7 */ (n141 ? (\pp[7]  ? n91 : !n91) : (\pp[7]  ? !n91 : n91));
assign n268 = /* LUT    7  3  3 */ n61;
assign n269 = /* LUT   11  1  5 */ (n139 ? (\pp[5]  ? n89 : !n89) : (\pp[5]  ? !n89 : n89));
assign n270 = /* LUT   11  1  3 */ (n137 ? (\pp[3]  ? n90 : !n90) : (\pp[3]  ? !n90 : n90));
assign n271 = /* LUT   11  2  3 */ (n146 ? (n103 ? \pp[11]  : !\pp[11] ) : (n103 ? !\pp[11]  : \pp[11] ));
assign n272 = /* LUT    6  3  6 */ (n38 ? (n60 ? (n34 ? n71 : 1'b0) : 1'b0) : 1'b0);
assign n273 = /* LUT   11  1  1 */ (n135 ? (n93 ? \pp[1]  : !\pp[1] ) : (n93 ? !\pp[1]  : \pp[1] ));
assign n274 = /* LUT   11  2  1 */ (n144 ? (\pp[9]  ? n106 : !n106) : (\pp[9]  ? !n106 : n106));
assign n275 = /* LUT   12  1  0 */ (\A[14]  ? (n134 ? 1'b1 : n1) : (n134 ? !n1 : 1'b0));
assign n276 = /* LUT    5  1  6 */ (n30 ? (\B[5]  ? 1'b1 : !n1) : (\B[5]  ? n1 : 1'b0));
assign n277 = /* LUT    9  2  3 */ (n79 ? (\B[8]  ? 1'b1 : !n1) : (\B[8]  ? n1 : 1'b0));
assign n278 = /* LUT   11  2  7 */ (n150 ? (n143 ? \pp[15]  : !\pp[15] ) : (n143 ? !\pp[15]  : \pp[15] ));
assign n279 = /* LUT    5  4  2 */ n59;
assign n280 = /* LUT    6  4  3 */ !n42;
assign n281 = /* LUT   11  2  5 */ (n148 ? (n134 ? \pp[13]  : !\pp[13] ) : (n134 ? !\pp[13]  : \pp[13] ));
assign n282 = /* LUT    5  4  0 */ (n47 ? 1'b0 : (n49 ? 1'b0 : n50));
assign n283 = /* LUT    5  1  2 */ (n29 ? (\B[4]  ? 1'b1 : !n1) : (\B[4]  ? n1 : 1'b0));
assign n284 = /* LUT    9  2  7 */ (n75 ? (\B[12]  ? 1'b1 : !n1) : (\B[12]  ? n1 : 1'b0));
assign n285 = /* LUT   11  4  4 */ (n178 ? (\pp[28]  ? n168 : !n168) : (\pp[28]  ? !n168 : n168));
assign n286 = /* LUT    5  4  6 */ (n57 ? 1'b1 : (n44 ? n56 : 1'b0));
assign n287 = /* LUT   12  3  7 */ n156;
assign n288 = /* LUT   11  4  6 */ (n180 ? (n22 ? n173 : !n173) : (n22 ? !n173 : n173));
assign n289 = /* LUT    5  4  4 */ !n59;
assign n290 = /* LUT   12  3  5 */ n152;
assign n291 = /* LUT   11  4  0 */ (n167 ? (\pp[24]  ? n170 : !n170) : (\pp[24]  ? !n170 : n170));
assign n292 = /* LUT   10  3  7 */ (\A[9]  ? (n1 ? 1'b1 : n104) : (n1 ? 1'b0 : n104));
assign n293 = /* LUT   12  3  3 */ n154;
assign n294 = /* LUT   11  3  0 */ (n151 ? (n156 ? \pp[16]  : !\pp[16] ) : (n156 ? !\pp[16]  : \pp[16] ));
assign n295 = /* LUT   11  4  2 */ (n176 ? (n169 ? \pp[26]  : !\pp[26] ) : (n169 ? !\pp[26]  : \pp[26] ));
assign n296 = /* LUT   10  3  1 */ (n103 ? (n1 ? \A[12]  : 1'b1) : (n1 ? \A[12]  : 1'b0));
assign n297 = /* LUT    5  2  5 */ (n53 ? (n1 ? \B[7]  : 1'b1) : (n1 ? \B[7]  : 1'b0));
assign n298 = /* LUT   12  3  1 */ n155;
assign n299 = /* LUT   11  3  2 */ (n161 ? (\pp[18]  ? n154 : !n154) : (\pp[18]  ? !n154 : n154));
assign n164 = /* CARRY 11  3  4 */ (\pp[20]  & n153) | ((\pp[20]  | n153) & n163);
assign n166 = /* CARRY 11  3  6 */ (\pp[22]  & n157) | ((\pp[22]  | n157) & n165);
assign n72  = /* CARRY  7  2  1 */ (1'b0 & n65) | ((1'b0 | n65) & n182);
assign n141 = /* CARRY 11  1  6 */ (n92 & \pp[6] ) | ((n92 | \pp[6] ) & n140);
assign n139 = /* CARRY 11  1  4 */ (\pp[4]  & n88) | ((\pp[4]  | n88) & n138);
assign n146 = /* CARRY 11  2  2 */ (n105 & \pp[10] ) | ((n105 | \pp[10] ) & n145);
assign n137 = /* CARRY 11  1  2 */ (\pp[2]  & n87) | ((\pp[2]  | n87) & n136);
assign n144 = /* CARRY 11  2  0 */ (\pp[8]  & n104) | ((\pp[8]  | n104) & n142);
assign n135 = /* CARRY 11  1  0 */ (n98 & \pp[0] ) | ((n98 | \pp[0] ) & n223);
assign n150 = /* CARRY 11  2  6 */ (\pp[14]  & n133) | ((\pp[14]  | n133) & n149);
assign n148 = /* CARRY 11  2  4 */ (n102 & \pp[12] ) | ((n102 | \pp[12] ) & n147);
assign n180 = /* CARRY 11  4  5 */ (\pp[29]  & n171) | ((\pp[29]  | n171) & n179);
assign n161 = /* CARRY 11  3  1 */ (n159 & \pp[17] ) | ((n159 | \pp[17] ) & n160);
assign n176 = /* CARRY 11  4  1 */ (\pp[25]  & n174) | ((\pp[25]  | n174) & n175);
assign n163 = /* CARRY 11  3  3 */ (\pp[19]  & n155) | ((\pp[19]  | n155) & n162);
assign n178 = /* CARRY 11  4  3 */ (\pp[27]  & n172) | ((\pp[27]  | n172) & n177);
assign n73  = /* CARRY  7  2  2 */ (1'b0 & n66) | ((1'b0 | n66) & n72);
assign n165 = /* CARRY 11  3  5 */ (n152 & \pp[21] ) | ((n152 | \pp[21] ) & n164);
assign n167 = /* CARRY 11  3  7 */ (n158 & \pp[23] ) | ((n158 | \pp[23] ) & n166);
assign n182 = /* CARRY  7  2  0 */ (1'b0 & n68) | ((1'b0 | n68) & n255);
assign n142 = /* CARRY 11  1  7 */ (n91 & \pp[7] ) | ((n91 | \pp[7] ) & n141);
assign n140 = /* CARRY 11  1  5 */ (n89 & \pp[5] ) | ((n89 | \pp[5] ) & n139);
assign n138 = /* CARRY 11  1  3 */ (n90 & \pp[3] ) | ((n90 | \pp[3] ) & n137);
assign n147 = /* CARRY 11  2  3 */ (\pp[11]  & n103) | ((\pp[11]  | n103) & n146);
assign n136 = /* CARRY 11  1  1 */ (\pp[1]  & n93) | ((\pp[1]  | n93) & n135);
assign n145 = /* CARRY 11  2  1 */ (n106 & \pp[9] ) | ((n106 | \pp[9] ) & n144);
assign n151 = /* CARRY 11  2  7 */ (\pp[15]  & n143) | ((\pp[15]  | n143) & n150);
assign n149 = /* CARRY 11  2  5 */ (\pp[13]  & n134) | ((\pp[13]  | n134) & n148);
assign n179 = /* CARRY 11  4  4 */ (n168 & \pp[28] ) | ((n168 | \pp[28] ) & n178);
assign n181 = /* CARRY 11  4  6 */ (n173 & n22) | ((n173 | n22) & n180);
assign n175 = /* CARRY 11  4  0 */ (n170 & \pp[24] ) | ((n170 | \pp[24] ) & n167);
assign n160 = /* CARRY 11  3  0 */ (\pp[16]  & n156) | ((\pp[16]  | n156) & n151);
assign n177 = /* CARRY 11  4  2 */ (\pp[26]  & n169) | ((\pp[26]  | n169) & n176);
assign n162 = /* CARRY 11  3  2 */ (n154 & \pp[18] ) | ((n154 | \pp[18] ) & n161);
/* FF 10  3  3 */ always @(negedge clk) if (n3) n103 <= 1'b0 ? 1'b0 : n183;
/* FF  5  2  7 */ always @(negedge clk) if (n3) n39 <= 1'b0 ? 1'b0 : n184;
/* FF  7  2  3 */ assign n63 = n185;
/* FF 11  3  4 */ always @(negedge clk) if (n2) \pp[20]  <= n1 ? 1'b0 : n186;
/* FF 10  1  6 */ always @(negedge clk) if (n3) n92 <= 1'b0 ? 1'b0 : n187;
/* FF  5  2  1 */ assign n34 = n188;
/* FF 11  3  6 */ always @(negedge clk) if (n2) \pp[22]  <= n1 ? 1'b0 : n189;
/* FF  7  2  1 */ assign n61 = n190;
/* FF 10  1  4 */ always @(negedge clk) if (n3) n90 <= 1'b0 ? 1'b0 : n191;
/* FF 10  1  2 */ always @(negedge clk) if (n3) n88 <= 1'b0 ? 1'b0 : n192;
/* FF 12  2  4 */ always @(negedge clk) if (n3) n143 <= 1'b0 ? 1'b0 : n193;
/* FF  9  1  1 */ always @(negedge clk) if (n3) n75 <= 1'b0 ? 1'b0 : n194;
/* FF  1 25  4 */ assign \pp[30]  = n195;
/* FF 12  4  6 */ always @(negedge clk) if (n3) n173 <= n1 ? 1'b0 : n196;
/* FF 10  1  0 */ always @(negedge clk) if (n3) n87 <= 1'b0 ? 1'b0 : n197;
/* FF  9  1  3 */ always @(negedge clk) if (n3) n76 <= 1'b0 ? 1'b0 : n198;
/* FF 12  4  4 */ always @(negedge clk) if (n3) n171 <= n1 ? 1'b0 : n199;
/* FF  7  3  4 */ always @(posedge clk) if (n64) n66 <= n27 ? 1'b0 : n200;
/* FF 10  2  6 */ always @(negedge clk) if (n3) n95 <= n99 ? 1'b0 : n201;
/* FF 12  4  2 */ always @(negedge clk) if (n3) n169 <= n1 ? 1'b0 : n202;
/* FF  7  3  6 */ always @(posedge clk) if (n64) n67 <= n27 ? 1'b0 : n203;
/* FF 10  2  4 */ assign n99 = n204;
/* FF  5  3  0 */ always @(posedge clk) if (n46) n40 <= 1'b0 ? 1'b0 : n205;
/* FF  6  3  1 */ always @(posedge clk) if (n59) n1 <= 1'b0 ? 1'b0 : n206;
/* FF  5  3  6 */ assign n42 = n207;
/* FF 11  1  6 */ always @(negedge clk) if (n2) \pp[6]  <= n1 ? 1'b0 : n208;
/* FF  7  3  2 */ assign n64 = n209;
/* FF  5  3  4 */ always @(posedge clk) if (n46) done <= 1'b0 ? 1'b0 : n210;
/* FF 11  1  4 */ always @(negedge clk) if (n2) \pp[4]  <= n1 ? 1'b0 : n211;
/* FF 11  2  2 */ always @(negedge clk) if (n2) \pp[10]  <= n1 ? 1'b0 : n212;
/* FF  6  3  5 */ always @(posedge clk) if (n59) n55 <= 1'b0 ? 1'b0 : n213;
/* FF 12  1  5 */ always @(negedge clk) if (n3) n134 <= 1'b0 ? 1'b0 : n214;
/* FF  9  2  0 */ always @(negedge clk) if (n3) n79 <= 1'b0 ? 1'b0 : n215;
/* FF  6  4  4 */ assign n59 = n216;
/* FF 11  1  2 */ always @(negedge clk) if (n2) \pp[2]  <= n1 ? 1'b0 : n217;
/* FF 11  2  0 */ always @(negedge clk) if (n2) \pp[8]  <= n1 ? 1'b0 : n218;
/* FF  6  3  7 */ assign n57 = n219;
/* FF  5  1  7 */ always @(negedge clk) if (n3) n30 <= 1'b0 ? 1'b0 : n220;
/* FF  9  2  2 */ assign n60 = n221;
/* FF 11  1  0 */ always @(negedge clk) if (n2) \pp[0]  <= n1 ? 1'b0 : n222;
/* FF 11  2  6 */ always @(negedge clk) if (n2) \pp[14]  <= n1 ? 1'b0 : n224;
/* FF  6  4  0 */ assign n58 = n225;
/* FF  9  2  4 */ always @(negedge clk) if (n3) n80 <= 1'b0 ? 1'b0 : n226;
/* FF 11  2  4 */ always @(negedge clk) if (n2) \pp[12]  <= n1 ? 1'b0 : n227;
/* FF  5  4  3 */ always @(posedge clk) if (1'b1) n47 <= n48 ? 1'b0 : n228;
/* FF  6  4  2 */ assign n2 = n229;
/* FF  9  2  6 */ always @(negedge clk) if (n3) n81 <= 1'b0 ? 1'b0 : n230;
/* FF  6  2  0 */ assign n3 = n231;
/* FF  5  4  1 */ assign n45 = n232;
/* FF 12  3  6 */ always @(negedge clk) if (n3) n158 <= n1 ? 1'b0 : n233;
/* FF 11  4  5 */ always @(negedge clk) if (n2) \pp[29]  <= n1 ? 1'b0 : n234;
/* FF 10  3  4 */ always @(negedge clk) if (n3) n104 <= 1'b0 ? 1'b0 : n235;
/* FF  5  4  7 */ always @(posedge clk) if (1'b1) n50 <= n48 ? 1'b0 : n236;
/* FF  9  3  3 */ assign n71 = n237;
/* FF 12  3  4 */ always @(negedge clk) if (n3) n156 <= n1 ? 1'b0 : n238;
/* FF 11  4  7 */ always @(negedge clk) if (n2) \pp[31]  <= n1 ? 1'b0 : n239;
/* FF 10  3  6 */ always @(negedge clk) if (n3) n105 <= 1'b0 ? 1'b0 : n240;
/* FF 12  3  2 */ always @(negedge clk) if (n3) n154 <= n1 ? 1'b0 : n241;
/* FF 11  3  1 */ always @(negedge clk) if (n2) \pp[17]  <= n1 ? 1'b0 : n242;
/* FF 11  4  1 */ always @(negedge clk) if (n2) \pp[25]  <= n1 ? 1'b0 : n243;
/* FF  5  2  4 */ always @(negedge clk) if (n3) n36 <= 1'b0 ? 1'b0 : n244;
/* FF 12  3  0 */ always @(negedge clk) if (n3) n152 <= n1 ? 1'b0 : n245;
/* FF 11  3  3 */ always @(negedge clk) if (n2) \pp[19]  <= n1 ? 1'b0 : n246;
/* FF 11  4  3 */ always @(negedge clk) if (n2) \pp[27]  <= n1 ? 1'b0 : n247;
/* FF  5  2  6 */ assign n38 = n248;
/* FF  7  2  2 */ assign n62 = n249;
/* FF 11  3  5 */ always @(negedge clk) if (n2) \pp[21]  <= n1 ? 1'b0 : n250;
/* FF  5  2  0 */ always @(negedge clk) if (n3) n33 <= 1'b0 ? 1'b0 : n251;
/* FF 11  3  7 */ always @(negedge clk) if (n2) \pp[23]  <= n1 ? 1'b0 : n252;
/* FF  7  2  0 */ assign n253 = n254;
/* FF 10  1  7 */ always @(negedge clk) if (n3) n93 <= 1'b0 ? 1'b0 : n256;
/* FF  5  2  2 */ always @(negedge clk) if (n3) n35 <= 1'b0 ? 1'b0 : n257;
/* FF 10  1  5 */ always @(negedge clk) if (n3) n91 <= 1'b0 ? 1'b0 : n258;
/* FF 12  4  7 */ always @(negedge clk) if (n3) n174 <= n1 ? 1'b0 : n259;
/* FF 10  1  3 */ always @(negedge clk) if (n3) n89 <= 1'b0 ? 1'b0 : n260;
/* FF 10  2  1 */ always @(negedge clk) if (n3) n98 <= n99 ? 1'b0 : n261;
/* FF 12  4  5 */ always @(negedge clk) if (n3) n172 <= n1 ? 1'b0 : n262;
/* FF 12  4  3 */ always @(negedge clk) if (n3) n170 <= n1 ? 1'b0 : n263;
/* FF  7  3  7 */ always @(posedge clk) if (n64) n68 <= n27 ? 1'b0 : n264;
/* FF 12  4  1 */ always @(negedge clk) if (n3) n168 <= n1 ? 1'b0 : n265;
/* FF  5  3  7 */ assign n43 = n266;
/* FF 11  1  7 */ always @(negedge clk) if (n2) \pp[7]  <= n1 ? 1'b0 : n267;
/* FF  7  3  3 */ always @(posedge clk) if (n64) n65 <= n27 ? 1'b0 : n268;
/* FF 11  1  5 */ always @(negedge clk) if (n2) \pp[5]  <= n1 ? 1'b0 : n269;
/* FF 11  1  3 */ always @(negedge clk) if (n2) \pp[3]  <= n1 ? 1'b0 : n270;
/* FF 11  2  3 */ always @(negedge clk) if (n2) \pp[11]  <= n1 ? 1'b0 : n271;
/* FF  6  3  6 */ assign n56 = n272;
/* FF 11  1  1 */ always @(negedge clk) if (n2) \pp[1]  <= n1 ? 1'b0 : n273;
/* FF 11  2  1 */ always @(negedge clk) if (n2) \pp[9]  <= n1 ? 1'b0 : n274;
/* FF 12  1  0 */ always @(negedge clk) if (n3) n133 <= 1'b0 ? 1'b0 : n275;
/* FF  5  1  6 */ always @(negedge clk) if (n3) n29 <= 1'b0 ? 1'b0 : n276;
/* FF  9  2  3 */ always @(negedge clk) if (n3) n53 <= 1'b0 ? 1'b0 : n277;
/* FF 11  2  7 */ always @(negedge clk) if (n2) \pp[15]  <= n1 ? 1'b0 : n278;
/* FF  5  4  2 */ assign n46 = n279;
/* FF  6  4  3 */ assign n27 = n280;
/* FF 11  2  5 */ always @(negedge clk) if (n2) \pp[13]  <= n1 ? 1'b0 : n281;
/* FF  5  4  0 */ assign n44 = n282;
/* FF  5  1  2 */ always @(negedge clk) if (n3) n28 <= 1'b0 ? 1'b0 : n283;
/* FF  9  2  7 */ always @(negedge clk) if (n3) n82 <= 1'b0 ? 1'b0 : n284;
/* FF 11  4  4 */ always @(negedge clk) if (n2) \pp[28]  <= n1 ? 1'b0 : n285;
/* FF  5  4  6 */ always @(posedge clk) if (1'b1) n49 <= n48 ? 1'b0 : n286;
/* FF 12  3  7 */ always @(negedge clk) if (n3) n159 <= n1 ? 1'b0 : n287;
/* FF 11  4  6 */ always @(negedge clk) if (n2) n22 <= n1 ? 1'b0 : n288;
/* FF  5  4  4 */ assign n48 = n289;
/* FF 12  3  5 */ always @(negedge clk) if (n3) n157 <= n1 ? 1'b0 : n290;
/* FF 11  4  0 */ always @(negedge clk) if (n2) \pp[24]  <= n1 ? 1'b0 : n291;
/* FF 10  3  7 */ always @(negedge clk) if (n3) n106 <= 1'b0 ? 1'b0 : n292;
/* FF 12  3  3 */ always @(negedge clk) if (n3) n155 <= n1 ? 1'b0 : n293;
/* FF 11  3  0 */ always @(negedge clk) if (n2) \pp[16]  <= n1 ? 1'b0 : n294;
/* FF 11  4  2 */ always @(negedge clk) if (n2) \pp[26]  <= n1 ? 1'b0 : n295;
/* FF 10  3  1 */ always @(negedge clk) if (n3) n102 <= 1'b0 ? 1'b0 : n296;
/* FF  5  2  5 */ always @(negedge clk) if (n3) n37 <= 1'b0 ? 1'b0 : n297;
/* FF 12  3  1 */ always @(negedge clk) if (n3) n153 <= n1 ? 1'b0 : n298;
/* FF 11  3  2 */ always @(negedge clk) if (n2) \pp[18]  <= n1 ? 1'b0 : n299;

endmodule

