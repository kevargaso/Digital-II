
//
// Verific Verilog Description of module SOC
//

module SOC (clk, resetn, LEDS, RXD, TXD);
    input clk /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input resetn /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output LEDS /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input RXD /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output TXD /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    
    
    wire n6, n7, n8, n9, \CPU/aluShamt[0] , \CPU/state[0] , n12, 
        n13, n14, n15, \RAM_rdata[24] , \CPU/rs1[16] , \CPU/rs1[17] , 
        \CPU/rs1[18] , \CPU/rs1[19] , \CPU/rs1[20] , \CPU/rs1[21] , 
        \CPU/rs1[22] , \CPU/rs1[23] , \CPU/rs1[24] , \CPU/rs1[25] , 
        \CPU/rs1[26] , \CPU/rs1[27] , \CPU/rs1[28] , \CPU/rs1[29] , 
        \CPU/rs1[30] , \CPU/rs1[31] , \CPU/rs1[0] , \CPU/rs1[1] , \CPU/rs1[2] , 
        \CPU/rs1[3] , \CPU/rs1[4] , \CPU/rs1[5] , \CPU/rs1[6] , \CPU/rs1[7] , 
        \CPU/rs1[8] , \CPU/rs1[9] , \CPU/rs1[10] , \CPU/rs1[11] , \CPU/rs1[12] , 
        \CPU/rs1[13] , \CPU/rs1[14] , \CPU/rs1[15] , \CPU/rs2[8] , \CPU/rs2[9] , 
        \CPU/rs2[10] , \CPU/rs2[11] , \CPU/rs2[12] , \CPU/rs2[13] , 
        \CPU/rs2[14] , \CPU/rs2[15] , \CPU/instr[2] , \CPU/cycles[0] , 
        \CPU/rs2[16] , \CPU/rs2[17] , \CPU/rs2[18] , \CPU/rs2[19] , 
        \CPU/rs2[20] , \CPU/rs2[21] , \CPU/rs2[22] , \CPU/rs2[23] , 
        \CPU/rs2[24] , \CPU/rs2[25] , \CPU/rs2[26] , \CPU/rs2[27] , 
        \CPU/rs2[28] , \CPU/rs2[29] , \CPU/rs2[30] , \CPU/rs2[31] , 
        \CPU/aluReg[1] , \CPU/aluReg[0] , \CPU/aluShamt[1] , \CPU/aluShamt[2] , 
        \CPU/aluShamt[3] , \CPU/aluShamt[4] , \CPU/state[1] , \CPU/state[2] , 
        \CPU/state[3] , \CPU/PC[1] , \CPU/PC[2] , \CPU/PC[3] , \CPU/PC[4] , 
        \CPU/PC[5] , \CPU/PC[6] , \CPU/PC[7] , \CPU/PC[8] , \CPU/PC[9] , 
        \CPU/PC[10] , \CPU/PC[11] , \CPU/PC[12] , \CPU/PC[13] , \CPU/PC[14] , 
        \CPU/PC[15] , \CPU/PC[16] , \CPU/PC[17] , \CPU/PC[18] , \CPU/PC[19] , 
        \CPU/PC[20] , \CPU/PC[21] , \CPU/PC[22] , \CPU/PC[23] , \CPU/instr[3] , 
        \CPU/instr[4] , \CPU/instr[5] , \CPU/instr[6] , \CPU/instr[7] , 
        \CPU/instr[8] , \CPU/instr[9] , \CPU/instr[10] , \CPU/instr[11] , 
        \CPU/instr[12] , \CPU/instr[13] , \CPU/instr[14] , \CPU/instr[15] , 
        \CPU/instr[16] , \CPU/instr[17] , \CPU/instr[18] , \CPU/instr[19] , 
        \CPU/instr[20] , \CPU/instr[21] , \CPU/instr[22] , \CPU/instr[23] , 
        \CPU/instr[24] , \CPU/instr[25] , \CPU/instr[26] , \CPU/instr[27] , 
        \CPU/instr[28] , \CPU/instr[29] , \CPU/instr[30] , \CPU/instr[31] , 
        \CPU/cycles[1] , \CPU/cycles[2] , \CPU/cycles[3] , \CPU/cycles[4] , 
        \CPU/cycles[5] , \CPU/cycles[6] , \CPU/cycles[7] , \CPU/cycles[8] , 
        \CPU/cycles[9] , \CPU/cycles[10] , \CPU/cycles[11] , \CPU/cycles[12] , 
        \CPU/cycles[13] , \CPU/cycles[14] , \CPU/cycles[15] , \CPU/cycles[16] , 
        \CPU/cycles[17] , \CPU/cycles[18] , \CPU/cycles[19] , \CPU/cycles[20] , 
        \CPU/cycles[21] , \CPU/cycles[22] , \CPU/cycles[23] , \CPU/cycles[24] , 
        \CPU/cycles[25] , \CPU/cycles[26] , \CPU/cycles[27] , \CPU/cycles[28] , 
        \CPU/cycles[29] , \CPU/cycles[30] , \CPU/cycles[31] , \CPU/aluReg[2] , 
        \CPU/aluReg[3] , \CPU/aluReg[4] , \CPU/aluReg[5] , \CPU/aluReg[6] , 
        \CPU/aluReg[7] , \CPU/aluReg[8] , \CPU/aluReg[9] , \CPU/aluReg[10] , 
        \CPU/aluReg[11] , \CPU/aluReg[12] , \CPU/aluReg[13] , \CPU/aluReg[14] , 
        \CPU/aluReg[15] , \CPU/aluReg[16] , \CPU/aluReg[17] , \CPU/aluReg[18] , 
        \CPU/aluReg[19] , \CPU/aluReg[20] , \CPU/aluReg[21] , \CPU/aluReg[22] , 
        \CPU/aluReg[23] , \CPU/aluReg[24] , \CPU/aluReg[25] , \CPU/aluReg[26] , 
        \CPU/aluReg[27] , \CPU/aluReg[28] , \CPU/aluReg[29] , \CPU/aluReg[30] , 
        \CPU/aluReg[31] , \RAM_rdata[2] , \RAM_rdata[16] , \RAM_rdata[25] , 
        \RAM_rdata[10] , n209, n210, \RAM_rdata[0] , \RAM_rdata[8] , 
        \RAM_rdata[26] , \RAM_rdata[18] , \RAM_rdata[27] , \RAM_rdata[28] , 
        \RAM_rdata[29] , \RAM_rdata[30] , \RAM_rdata[31] , \RAM_rdata[17] , 
        \RAM_rdata[19] , \RAM_rdata[20] , \RAM_rdata[21] , \RAM_rdata[22] , 
        \RAM_rdata[23] , \RAM_rdata[9] , \RAM_rdata[11] , \RAM_rdata[12] , 
        \RAM_rdata[13] , \RAM_rdata[14] , \RAM_rdata[15] , \RAM_rdata[1] , 
        \RAM_rdata[3] , \RAM_rdata[4] , \RAM_rdata[5] , \RAM_rdata[6] , 
        \RAM_rdata[7] , n238, n239, \per_uart/uart_ctrl[0] , \uart_dout[0] , 
        \per_uart/d_in_uart[0] , \per_uart/uart_ctrl[1] , \uart_dout[1] , 
        \uart_dout[2] , \uart_dout[3] , \uart_dout[4] , \uart_dout[5] , 
        \uart_dout[6] , \uart_dout[7] , \uart_dout[8] , \uart_dout[9] , 
        \per_uart/uart0/uart_rxd1 , \per_uart/uart0/uart_rxd2 , \per_uart/uart0/rx_busy , 
        \per_uart/uart0/rx_count16[0] , \per_uart/uart0/rx_bitcount[0] , 
        \per_uart/rx_data[0] , \per_uart/rx_avail , \per_uart/rx_error , 
        \per_uart/tx_busy , \per_uart/uart0/tx_count16[0] , \per_uart/uart0/txd_reg[0] , 
        \per_uart/uart0/tx_bitcount[0] , \per_uart/uart0/enable16_counter[0] , 
        \per_uart/uart0/rx_count16[1] , \per_uart/uart0/rx_count16[2] , 
        \per_uart/uart0/rx_count16[3] , \per_uart/uart0/rx_bitcount[1] , 
        \per_uart/uart0/rx_bitcount[2] , \per_uart/uart0/rx_bitcount[3] , 
        \per_uart/rx_data[1] , \per_uart/rx_data[2] , \per_uart/rx_data[3] , 
        \per_uart/rx_data[4] , \per_uart/rx_data[5] , \per_uart/rx_data[6] , 
        \per_uart/rx_data[7] , \per_uart/uart0/tx_count16[1] , \per_uart/uart0/tx_count16[2] , 
        \per_uart/uart0/tx_count16[3] , \per_uart/uart0/txd_reg[1] , \per_uart/uart0/txd_reg[2] , 
        \per_uart/uart0/txd_reg[3] , \per_uart/uart0/txd_reg[4] , \per_uart/uart0/txd_reg[5] , 
        \per_uart/uart0/txd_reg[6] , \per_uart/uart0/txd_reg[7] , \per_uart/uart0/tx_bitcount[1] , 
        \per_uart/uart0/tx_bitcount[2] , \per_uart/uart0/tx_bitcount[3] , 
        \per_uart/uart0/enable16_counter[1] , \per_uart/uart0/enable16_counter[2] , 
        \per_uart/uart0/enable16_counter[3] , \per_uart/uart0/enable16_counter[4] , 
        \per_uart/d_in_uart[1] , \per_uart/d_in_uart[2] , \per_uart/d_in_uart[3] , 
        \per_uart/d_in_uart[4] , \per_uart/d_in_uart[5] , \per_uart/d_in_uart[6] , 
        \per_uart/d_in_uart[7] , \mult1/A[0] , \mult1/B[0] , \mult_dout[0] , 
        \mult1/init , \mult1/A[1] , \mult1/A[2] , \mult1/A[3] , \mult1/A[4] , 
        \mult1/A[5] , \mult1/A[6] , \mult1/A[7] , \mult1/A[8] , \mult1/A[9] , 
        \mult1/A[10] , \mult1/A[11] , \mult1/A[12] , \mult1/A[13] , 
        \mult1/A[14] , \mult1/A[15] , \mult1/B[1] , \mult1/B[2] , \mult1/B[3] , 
        \mult1/B[4] , \mult1/B[5] , \mult1/B[6] , \mult1/B[7] , \mult1/B[8] , 
        \mult1/B[9] , \mult1/B[10] , \mult1/B[11] , \mult1/B[12] , \mult1/B[13] , 
        \mult1/B[14] , \mult1/B[15] , \mult_dout[1] , \mult_dout[2] , 
        \mult_dout[3] , \mult_dout[4] , \mult_dout[5] , \mult_dout[6] , 
        \mult_dout[7] , \mult_dout[8] , \mult_dout[9] , \mult_dout[10] , 
        \mult_dout[11] , \mult_dout[12] , \mult_dout[13] , \mult_dout[14] , 
        \mult_dout[15] , \mult_dout[16] , \mult_dout[17] , \mult_dout[18] , 
        \mult_dout[19] , \mult_dout[20] , \mult_dout[21] , \mult_dout[22] , 
        \mult_dout[23] , \mult_dout[24] , \mult_dout[25] , \mult_dout[26] , 
        \mult_dout[27] , \mult_dout[28] , \mult_dout[29] , \mult_dout[30] , 
        \mult_dout[31] , \mult1/result[0] , \mult1/mult1/state[0] , \mult1/mult1/A[0] , 
        \mult1/mult1/B[0] , \mult1/mult1/count[0] , \mult1/done , \mult1/result[1] , 
        \mult1/result[2] , \mult1/result[3] , \mult1/result[4] , \mult1/result[5] , 
        \mult1/result[6] , \mult1/result[7] , \mult1/result[8] , \mult1/result[9] , 
        \mult1/result[10] , \mult1/result[11] , \mult1/result[12] , \mult1/result[13] , 
        \mult1/result[14] , \mult1/result[15] , \mult1/result[16] , \mult1/result[17] , 
        \mult1/result[18] , \mult1/result[19] , \mult1/result[20] , \mult1/result[21] , 
        \mult1/result[22] , \mult1/result[23] , \mult1/result[24] , \mult1/result[25] , 
        \mult1/result[26] , \mult1/result[27] , \mult1/result[28] , \mult1/result[29] , 
        \mult1/result[30] , \mult1/result[31] , \mult1/mult1/state[1] , 
        \mult1/mult1/state[2] , \mult1/mult1/A[1] , \mult1/mult1/A[2] , 
        \mult1/mult1/A[3] , \mult1/mult1/A[4] , \mult1/mult1/A[5] , \mult1/mult1/A[6] , 
        \mult1/mult1/A[7] , \mult1/mult1/A[8] , \mult1/mult1/A[9] , \mult1/mult1/A[10] , 
        \mult1/mult1/A[11] , \mult1/mult1/A[12] , \mult1/mult1/A[13] , 
        \mult1/mult1/A[14] , \mult1/mult1/A[15] , \mult1/mult1/B[1] , 
        \mult1/mult1/B[2] , \mult1/mult1/B[3] , \mult1/mult1/B[4] , \mult1/mult1/B[5] , 
        \mult1/mult1/B[6] , \mult1/mult1/B[7] , \mult1/mult1/B[8] , \mult1/mult1/B[9] , 
        \mult1/mult1/B[10] , \mult1/mult1/B[11] , \mult1/mult1/B[12] , 
        \mult1/mult1/B[13] , \mult1/mult1/B[14] , \mult1/mult1/B[15] , 
        \mult1/mult1/count[1] , \mult1/mult1/count[2] , \mult1/mult1/count[3] , 
        \mult1/mult1/count[4] , n451, n452, n453, n454, n455, n456, 
        n457, n458, n459, n460, n461, n462, n463, n464, n465, 
        n466, n467, n468, n469, n470, n471, n472, n473, n474, 
        n475, n476, n477, n478, n479, n480, n481, n482, n483, 
        n484, n485, n486, n487, n488, n489, n490, n491, n492, 
        n493, n494, n495, n496, n497, n498, n499, n500, n501, 
        n502, n503, n504, n505, n506, n507, n508, n509, n510, 
        n511, n512, n513, n514, n515, n516, n517, n518, n519, 
        n520, n521, n522, n523, n524, n525, n526, n527, n528, 
        n529, n530, n531, n532, n533, n534, n535, n536, n537, 
        n538, n539, n540, n541, n542, n543, n544, n545, n546, 
        n547, n548, n549, n550, n551, n552, n553, n554, n555, 
        n556, n557, n558, n559, n560, n561, n562, n563, n564, 
        n565, n566, n567, n568, n569, n570, n571, n572, n573, 
        n574, n575, n576, n577, n578, n579, n580, n581, n582, 
        n583, n584, n585, n586, n587, n588, n589, n590, n591, 
        n592, n593, n594, n595, n596, n597, n598, n599, n600, 
        n601, n602, n603, n604, n605, n606, n607, n608, n609, 
        n610, n611, n612, n613, n614, n615, n616, n617, n618, 
        n619, n620, n621, n622, n623, n624, n625, n626, n627, 
        n628, n629, n630, n631, n632, n633, n634, n635, n636, 
        n637, n638, n639, n640, n641, n642, n643, n644, n645, 
        n646, n647, n648, n649, n650, n651, n652, n653, n654, 
        n655, n656, n657, n658, n659, n660, n661, n662, n663, 
        n664, n665, n666, n667, n668, n669, n670, n671, n672, 
        n673, n674, n675, n676, n677, n678, n679, n680, n681, 
        n682, n683, n684, n685, n686, n687, n688, n689, n690, 
        n691, n692, n693, n694, n695, n696, n697, n698, n699, 
        n700, n701, n702, n703, n704, n705, n706, n707, n708, 
        n709, n710, n711, n712, n713, n714, n715, n716, n717, 
        n718, n719, n720, n721, n722, n723, n724, n725, n726, 
        n727, n728, n729, n730, n731, n732, n733, n734, n735, 
        n736, n737, n738, n739, n740, n741, n742, n743, n744, 
        n745, n746, n747, n748, n749, n750, n751, n752, n753, 
        n754, n755, n756, n757, n758, n759, n760, n761, n762, 
        n763, n764, n765, n766, n767, n768, n769, n770, n771, 
        n772, n773, n774, n775, n776, n777, n778, n779, n780, 
        n781, n787, \CPU/n1034 , ceg_net77, \CPU/n2185 , n793, n107, 
        \mem_addr[2] , \mem_addr[3] , \mem_addr[4] , \mem_addr[5] , 
        \mem_addr[6] , \mem_addr[7] , \mem_addr[8] , \mem_addr[9] , 
        \mem_addr[10] , \mem_addr[11] , \mem_addr[12] , \mem_addr[13] , 
        \mem_wdata[24] , \RAM/n116 , \CPU/n3447 , \mem_rdata[15] , \mem_rdata[16] , 
        \mem_rdata[17] , \mem_rdata[18] , \mem_rdata[19] , \CPU/writeBackData[16] , 
        \CPU/writeBackData[17] , \CPU/writeBackData[18] , \CPU/writeBackData[19] , 
        \CPU/writeBackData[20] , \CPU/writeBackData[21] , \CPU/writeBackData[22] , 
        \CPU/writeBackData[23] , \CPU/writeBackData[24] , \CPU/writeBackData[25] , 
        \CPU/writeBackData[26] , \CPU/writeBackData[27] , \CPU/writeBackData[28] , 
        \CPU/writeBackData[29] , \CPU/writeBackData[30] , \CPU/writeBackData[31] , 
        \CPU/not_equal_22/n9 , \CPU/writeBack , \CPU/writeBackData[0] , 
        \CPU/writeBackData[1] , \CPU/writeBackData[2] , \CPU/writeBackData[3] , 
        \CPU/writeBackData[4] , \CPU/writeBackData[5] , \CPU/writeBackData[6] , 
        \CPU/writeBackData[7] , \CPU/writeBackData[8] , \CPU/writeBackData[9] , 
        \CPU/writeBackData[10] , \CPU/writeBackData[11] , \CPU/writeBackData[12] , 
        \CPU/writeBackData[13] , \CPU/writeBackData[14] , \CPU/writeBackData[15] , 
        \mem_rdata[20] , \mem_rdata[21] , \mem_rdata[22] , \mem_rdata[23] , 
        \mem_rdata[24] , \mem_rdata[2] , \CPU/n1066 , \CPU/n1067 , \CPU/n1033 , 
        \CPU/n1032 , \CPU/n1031 , \CPU/n1030 , \CPU/select_174/Select_1/n5 , 
        \CPU/n2183 , \CPU/n2182 , \CPU/n2063 , ceg_net32, \CPU/n2062 , 
        \CPU/n2061 , \CPU/n2060 , \CPU/n2059 , \CPU/n2058 , \CPU/n2057 , 
        \CPU/n2056 , \CPU/n2055 , \CPU/n2054 , \CPU/n2053 , \CPU/n2052 , 
        \CPU/n2051 , \CPU/n2050 , \CPU/n2049 , \CPU/n2048 , \CPU/n2047 , 
        \CPU/n2046 , \CPU/n2045 , \CPU/n2044 , \CPU/n2043 , \CPU/n2042 , 
        \CPU/n2041 , \mem_rdata[3] , \mem_rdata[4] , \mem_rdata[5] , 
        \mem_rdata[6] , \mem_rdata[7] , \mem_rdata[8] , \mem_rdata[9] , 
        \mem_rdata[10] , \mem_rdata[11] , \mem_rdata[12] , \mem_rdata[13] , 
        \mem_rdata[14] , \mem_rdata[25] , \mem_rdata[26] , \mem_rdata[27] , 
        \mem_rdata[28] , \mem_rdata[29] , \mem_rdata[30] , \mem_rdata[31] , 
        \CPU/n1065 , \CPU/n1064 , \CPU/n1063 , \CPU/n1062 , \CPU/n1061 , 
        \CPU/n1060 , \CPU/n1059 , \CPU/n1058 , \CPU/n1057 , \CPU/n1056 , 
        \CPU/n1055 , \CPU/n1054 , \CPU/n1053 , \CPU/n1052 , \CPU/n1051 , 
        \CPU/n1050 , \CPU/n1049 , \CPU/n1048 , \CPU/n1047 , \CPU/n1046 , 
        \CPU/n1045 , \CPU/n1044 , \CPU/n1043 , \CPU/n1042 , \CPU/n1041 , 
        \CPU/n1040 , \CPU/n1039 , \CPU/n1038 , \CPU/n1037 , \CPU/n1036 , 
        \mem_wdata[2] , \RAM/n104 , \mem_wdata[16] , \RAM/n112 , \mem_wdata[25] , 
        \mem_wdata[10] , \RAM/n108 , \mem_wdata[0] , \mem_wdata[8] , 
        \mem_wdata[26] , \mem_wdata[18] , \mem_wdata[27] , \mem_wdata[28] , 
        \mem_wdata[29] , \mem_wdata[30] , \mem_wdata[31] , \mem_wdata[17] , 
        \mem_wdata[19] , \mem_wdata[20] , \mem_wdata[21] , \mem_wdata[22] , 
        \mem_wdata[23] , \mem_wdata[9] , \mem_wdata[11] , \mem_wdata[12] , 
        \mem_wdata[13] , \mem_wdata[14] , \mem_wdata[15] , \mem_wdata[1] , 
        \mem_wdata[3] , \mem_wdata[4] , \mem_wdata[5] , \mem_wdata[6] , 
        \mem_wdata[7] , \per_uart/n25 , \per_uart/select_21/Select_0/n3 , 
        \per_uart/n15 , \per_uart/select_21/Select_1/n3 , \per_uart/select_21/Select_2/n3 , 
        \per_uart/select_21/Select_3/n3 , \per_uart/select_21/Select_4/n3 , 
        \per_uart/select_21/Select_5/n3 , \per_uart/select_21/Select_6/n3 , 
        \per_uart/select_21/Select_7/n4 , \per_uart/select_21/Select_8/n2 , 
        \per_uart/select_21/Select_9/n2 , \per_uart/uart0/n190 , ceg_net530, 
        \per_uart/uart0/n195 , ceg_net176, \per_uart/uart0/n200 , \per_uart/uart0/rxd_reg[0] , 
        \per_uart/uart0/n581 , \per_uart/uart0/n576 , ceg_net140, \per_uart/uart0/n242 , 
        ceg_net144, \per_uart/uart0/rxd_reg[1] , \per_uart/uart0/n582 , 
        \per_uart/uart0/n316 , \per_uart/uart0/n601 , \per_uart/uart0/n422 , 
        ceg_net203, \per_uart/uart0/n386 , ceg_net155, \per_uart/uart0/n438 , 
        ceg_net159, \per_uart/uart0/n427 , ceg_net246, \per_uart/uart0/n552 , 
        \per_uart/uart0/n194 , \per_uart/uart0/n193 , \per_uart/uart0/n192 , 
        \per_uart/uart0/n199 , \per_uart/uart0/n198 , \per_uart/uart0/n197 , 
        \per_uart/uart0/rxd_reg[2] , \per_uart/uart0/rxd_reg[3] , \per_uart/uart0/rxd_reg[4] , 
        \per_uart/uart0/rxd_reg[5] , \per_uart/uart0/rxd_reg[6] , \per_uart/uart0/rxd_reg[7] , 
        \per_uart/uart0/n421 , \per_uart/uart0/n420 , \per_uart/uart0/n419 , 
        \per_uart/uart0/n437 , \per_uart/uart0/n436 , \per_uart/uart0/n435 , 
        \per_uart/uart0/n434 , \per_uart/uart0/n433 , \per_uart/uart0/n432 , 
        \per_uart/uart0/n431 , \per_uart/uart0/n426 , \per_uart/uart0/n425 , 
        \per_uart/uart0/n424 , \per_uart/uart0/n732 , \per_uart/uart0/n737 , 
        \per_uart/uart0/n742 , \per_uart/uart0/n747 , \mult1/n402 , \mult1/n403 , 
        \mult1/n201 , \mult1/n165 , \mult1/n404 , \mult1/n200 , \mult1/n199 , 
        \mult1/n198 , \mult1/n197 , \mult1/n196 , \mult1/n195 , \mult1/n194 , 
        \mult1/n193 , \mult1/n192 , \mult1/n191 , \mult1/n190 , \mult1/n189 , 
        \mult1/n188 , \mult1/n187 , \mult1/n186 , \mult1/n185 , \mult1/n184 , 
        \mult1/n183 , \mult1/n182 , \mult1/n181 , \mult1/n180 , \mult1/n179 , 
        \mult1/n178 , \mult1/n177 , \mult1/n176 , \mult1/n175 , \mult1/n174 , 
        \mult1/n173 , \mult1/n172 , \mult1/n171 , \mult1/n170 , \mult1/mult1/n132 , 
        ceg_net913, \mult1/mult1/n64 , ceg_net252, \mult1/mult1/n81 , 
        ceg_net839, \mult1/mult1/n98 , \mult1/mult1/n138 , ceg_net847, 
        \mult1/mult1/n99 , ceg_net564, \mult1/mult1/n131 , \mult1/mult1/n130 , 
        \mult1/mult1/n129 , \mult1/mult1/n128 , \mult1/mult1/n127 , \mult1/mult1/n126 , 
        \mult1/mult1/n125 , \mult1/mult1/n124 , \mult1/mult1/n123 , \mult1/mult1/n122 , 
        \mult1/mult1/n121 , \mult1/mult1/n120 , \mult1/mult1/n119 , \mult1/mult1/n118 , 
        \mult1/mult1/n117 , \mult1/mult1/n116 , \mult1/mult1/n115 , \mult1/mult1/n114 , 
        \mult1/mult1/n113 , \mult1/mult1/n112 , \mult1/mult1/n111 , \mult1/mult1/n110 , 
        \mult1/mult1/n109 , \mult1/mult1/n108 , \mult1/mult1/n107 , \mult1/mult1/n106 , 
        \mult1/mult1/n105 , \mult1/mult1/n104 , \mult1/mult1/n103 , \mult1/mult1/n102 , 
        \mult1/mult1/n101 , \mult1/mult1/n63 , \mult1/mult1/n62 , \mult1/mult1/n80 , 
        \mult1/mult1/n79 , \mult1/mult1/n78 , \mult1/mult1/n77 , \mult1/mult1/n76 , 
        \mult1/mult1/n75 , \mult1/mult1/n74 , \mult1/mult1/n73 , \mult1/mult1/n72 , 
        \mult1/mult1/n71 , \mult1/mult1/n70 , \mult1/mult1/n69 , \mult1/mult1/n68 , 
        \mult1/mult1/n67 , \mult1/mult1/n66 , \mult1/mult1/n97 , \mult1/mult1/n96 , 
        \mult1/mult1/n95 , \mult1/mult1/n94 , \mult1/mult1/n93 , \mult1/mult1/n92 , 
        \mult1/mult1/n91 , \mult1/mult1/n90 , \mult1/mult1/n89 , \mult1/mult1/n88 , 
        \mult1/mult1/n87 , \mult1/mult1/n86 , \mult1/mult1/n85 , \mult1/mult1/n84 , 
        \mult1/mult1/n83 , \mult1/mult1/n137 , \mult1/mult1/n136 , \mult1/mult1/n135 , 
        \mult1/mult1/n134 , n1378, n1381, n1384, n1387, n1390, n1393, 
        n1396, n1399, n1402, n1405, n1408, n1411, n1414, n1417, 
        n1420, n1423, n1426, n1429, n1432, n1435, n1438, n1441, 
        n1444, n1447, n1450, n1453, n1525, n1527, n1529, n1531, 
        n1533, n1535, n1537, n1539, n1541, n1543, n1545, n1547, 
        n1549, n1551, n1553, n1555, n1557, n1559, n1561, n1563, 
        n1565, n1567, n1569, n1571, n1573, n1575, n1577, \clk~O , 
        n1579, n2159, n1581, \CPU/instr[4]~FF_frt_1_frt_2_q , n1583, 
        \CPU/instr[4]~FF_frt_1_q , n1585, \CPU/instr[2]~FF_frt_0_q , n1587, 
        n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, 
        n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, 
        n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, 
        n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, 
        n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, 
        n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, 
        n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, 
        n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, 
        n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, 
        n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, 
        n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, 
        n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, 
        n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, 
        n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, 
        n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, 
        n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, 
        n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, 
        n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, 
        n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, 
        n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, 
        n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, 
        n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, 
        n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, 
        n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, 
        n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, 
        n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, 
        n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, 
        n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, 
        n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, 
        n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, 
        n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, 
        n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, 
        n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, 
        n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, 
        n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, 
        n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, 
        n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, 
        n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, 
        n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, 
        n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, 
        n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, 
        n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, 
        n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, 
        n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, 
        n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, 
        n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, 
        n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, 
        n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, 
        n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, 
        n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, 
        n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, 
        n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, 
        n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, 
        n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, 
        n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, 
        n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, 
        n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, 
        n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, 
        n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, 
        n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, 
        n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, 
        n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, 
        n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, 
        n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, 
        n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, 
        n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, 
        n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, 
        n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, 
        n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, 
        n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, 
        n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, 
        n2157, n2158;
    
    EFX_FF \CPU/aluShamt[0]~FF  (.D(\CPU/n1034 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluShamt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluShamt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluShamt[0]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluShamt[0]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluShamt[0]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluShamt[0]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluShamt[0]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluShamt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/state[0]~FF  (.D(\CPU/n2185 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(resetn), .Q(\CPU/state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/state[0]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/state[0]~FF .SR_POLARITY = 1'b0;
    defparam \CPU/state[0]~FF .D_POLARITY = 1'b1;
    defparam \CPU/state[0]~FF .SR_SYNC = 1'b1;
    defparam \CPU/state[0]~FF .SR_VALUE = 1'b0;
    defparam \CPU/state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/instr[2]~FF  (.D(\mem_rdata[2] ), .CE(\CPU/n3447 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/instr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/instr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/instr[2]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/instr[2]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/instr[2]~FF .D_POLARITY = 1'b1;
    defparam \CPU/instr[2]~FF .SR_SYNC = 1'b1;
    defparam \CPU/instr[2]~FF .SR_VALUE = 1'b0;
    defparam \CPU/instr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/cycles[0]~FF  (.D(\CPU/cycles[0] ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/cycles[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/cycles[0]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/cycles[0]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/cycles[0]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/cycles[0]~FF .D_POLARITY = 1'b0;
    defparam \CPU/cycles[0]~FF .SR_SYNC = 1'b1;
    defparam \CPU/cycles[0]~FF .SR_VALUE = 1'b0;
    defparam \CPU/cycles[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/aluReg[1]~FF  (.D(\CPU/n1066 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluReg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluReg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluReg[1]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluReg[1]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluReg[1]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluReg[1]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluReg[1]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluReg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/aluReg[0]~FF  (.D(\CPU/n1067 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluReg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluReg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluReg[0]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluReg[0]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluReg[0]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluReg[0]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluReg[0]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluReg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/aluShamt[1]~FF  (.D(\CPU/n1033 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluShamt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluShamt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluShamt[1]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluShamt[1]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluShamt[1]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluShamt[1]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluShamt[1]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluShamt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/aluShamt[2]~FF  (.D(\CPU/n1032 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluShamt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluShamt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluShamt[2]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluShamt[2]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluShamt[2]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluShamt[2]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluShamt[2]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluShamt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/aluShamt[3]~FF  (.D(\CPU/n1031 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluShamt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluShamt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluShamt[3]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluShamt[3]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluShamt[3]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluShamt[3]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluShamt[3]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluShamt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/aluShamt[4]~FF  (.D(\CPU/n1030 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluShamt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluShamt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluShamt[4]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluShamt[4]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluShamt[4]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluShamt[4]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluShamt[4]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluShamt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/state[1]~FF  (.D(\CPU/select_174/Select_1/n5 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(resetn), .Q(\CPU/state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/state[1]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/state[1]~FF .SR_POLARITY = 1'b0;
    defparam \CPU/state[1]~FF .D_POLARITY = 1'b1;
    defparam \CPU/state[1]~FF .SR_SYNC = 1'b1;
    defparam \CPU/state[1]~FF .SR_VALUE = 1'b0;
    defparam \CPU/state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/state[2]~FF  (.D(\CPU/n2183 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(resetn), .Q(\CPU/state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/state[2]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/state[2]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/state[2]~FF .SR_POLARITY = 1'b0;
    defparam \CPU/state[2]~FF .D_POLARITY = 1'b1;
    defparam \CPU/state[2]~FF .SR_SYNC = 1'b1;
    defparam \CPU/state[2]~FF .SR_VALUE = 1'b0;
    defparam \CPU/state[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/state[3]~FF  (.D(\CPU/n2182 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(resetn), .Q(\CPU/state[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/state[3]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/state[3]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/state[3]~FF .SR_POLARITY = 1'b0;
    defparam \CPU/state[3]~FF .D_POLARITY = 1'b1;
    defparam \CPU/state[3]~FF .SR_SYNC = 1'b1;
    defparam \CPU/state[3]~FF .SR_VALUE = 1'b1;
    defparam \CPU/state[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/PC[1]~FF  (.D(\CPU/n2063 ), .CE(ceg_net32), .CLK(\clk~O ), 
           .SR(resetn), .Q(\CPU/PC[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/PC[1]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/PC[1]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/PC[1]~FF .SR_POLARITY = 1'b0;
    defparam \CPU/PC[1]~FF .D_POLARITY = 1'b1;
    defparam \CPU/PC[1]~FF .SR_SYNC = 1'b1;
    defparam \CPU/PC[1]~FF .SR_VALUE = 1'b0;
    defparam \CPU/PC[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/PC[2]~FF  (.D(\CPU/n2062 ), .CE(\CPU/state[2] ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\CPU/PC[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/PC[2]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/PC[2]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/PC[2]~FF .SR_POLARITY = 1'b0;
    defparam \CPU/PC[2]~FF .D_POLARITY = 1'b1;
    defparam \CPU/PC[2]~FF .SR_SYNC = 1'b1;
    defparam \CPU/PC[2]~FF .SR_VALUE = 1'b0;
    defparam \CPU/PC[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/PC[3]~FF  (.D(\CPU/n2061 ), .CE(\CPU/state[2] ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\CPU/PC[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/PC[3]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/PC[3]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/PC[3]~FF .SR_POLARITY = 1'b0;
    defparam \CPU/PC[3]~FF .D_POLARITY = 1'b1;
    defparam \CPU/PC[3]~FF .SR_SYNC = 1'b1;
    defparam \CPU/PC[3]~FF .SR_VALUE = 1'b0;
    defparam \CPU/PC[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/PC[4]~FF  (.D(\CPU/n2060 ), .CE(\CPU/state[2] ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\CPU/PC[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/PC[4]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/PC[4]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/PC[4]~FF .SR_POLARITY = 1'b0;
    defparam \CPU/PC[4]~FF .D_POLARITY = 1'b1;
    defparam \CPU/PC[4]~FF .SR_SYNC = 1'b1;
    defparam \CPU/PC[4]~FF .SR_VALUE = 1'b0;
    defparam \CPU/PC[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/PC[5]~FF  (.D(\CPU/n2059 ), .CE(\CPU/state[2] ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\CPU/PC[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/PC[5]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/PC[5]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/PC[5]~FF .SR_POLARITY = 1'b0;
    defparam \CPU/PC[5]~FF .D_POLARITY = 1'b1;
    defparam \CPU/PC[5]~FF .SR_SYNC = 1'b1;
    defparam \CPU/PC[5]~FF .SR_VALUE = 1'b0;
    defparam \CPU/PC[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/PC[6]~FF  (.D(\CPU/n2058 ), .CE(\CPU/state[2] ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\CPU/PC[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/PC[6]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/PC[6]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/PC[6]~FF .SR_POLARITY = 1'b0;
    defparam \CPU/PC[6]~FF .D_POLARITY = 1'b1;
    defparam \CPU/PC[6]~FF .SR_SYNC = 1'b1;
    defparam \CPU/PC[6]~FF .SR_VALUE = 1'b0;
    defparam \CPU/PC[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/PC[7]~FF  (.D(\CPU/n2057 ), .CE(\CPU/state[2] ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\CPU/PC[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/PC[7]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/PC[7]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/PC[7]~FF .SR_POLARITY = 1'b0;
    defparam \CPU/PC[7]~FF .D_POLARITY = 1'b1;
    defparam \CPU/PC[7]~FF .SR_SYNC = 1'b1;
    defparam \CPU/PC[7]~FF .SR_VALUE = 1'b0;
    defparam \CPU/PC[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/PC[8]~FF  (.D(\CPU/n2056 ), .CE(\CPU/state[2] ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\CPU/PC[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/PC[8]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/PC[8]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/PC[8]~FF .SR_POLARITY = 1'b0;
    defparam \CPU/PC[8]~FF .D_POLARITY = 1'b1;
    defparam \CPU/PC[8]~FF .SR_SYNC = 1'b1;
    defparam \CPU/PC[8]~FF .SR_VALUE = 1'b0;
    defparam \CPU/PC[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/PC[9]~FF  (.D(\CPU/n2055 ), .CE(\CPU/state[2] ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\CPU/PC[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/PC[9]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/PC[9]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/PC[9]~FF .SR_POLARITY = 1'b0;
    defparam \CPU/PC[9]~FF .D_POLARITY = 1'b1;
    defparam \CPU/PC[9]~FF .SR_SYNC = 1'b1;
    defparam \CPU/PC[9]~FF .SR_VALUE = 1'b0;
    defparam \CPU/PC[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/PC[10]~FF  (.D(\CPU/n2054 ), .CE(\CPU/state[2] ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\CPU/PC[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/PC[10]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/PC[10]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/PC[10]~FF .SR_POLARITY = 1'b0;
    defparam \CPU/PC[10]~FF .D_POLARITY = 1'b1;
    defparam \CPU/PC[10]~FF .SR_SYNC = 1'b1;
    defparam \CPU/PC[10]~FF .SR_VALUE = 1'b0;
    defparam \CPU/PC[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/PC[11]~FF  (.D(\CPU/n2053 ), .CE(\CPU/state[2] ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\CPU/PC[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/PC[11]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/PC[11]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/PC[11]~FF .SR_POLARITY = 1'b0;
    defparam \CPU/PC[11]~FF .D_POLARITY = 1'b1;
    defparam \CPU/PC[11]~FF .SR_SYNC = 1'b1;
    defparam \CPU/PC[11]~FF .SR_VALUE = 1'b0;
    defparam \CPU/PC[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/PC[12]~FF  (.D(\CPU/n2052 ), .CE(\CPU/state[2] ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\CPU/PC[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/PC[12]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/PC[12]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/PC[12]~FF .SR_POLARITY = 1'b0;
    defparam \CPU/PC[12]~FF .D_POLARITY = 1'b1;
    defparam \CPU/PC[12]~FF .SR_SYNC = 1'b1;
    defparam \CPU/PC[12]~FF .SR_VALUE = 1'b0;
    defparam \CPU/PC[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/PC[13]~FF  (.D(\CPU/n2051 ), .CE(\CPU/state[2] ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\CPU/PC[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/PC[13]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/PC[13]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/PC[13]~FF .SR_POLARITY = 1'b0;
    defparam \CPU/PC[13]~FF .D_POLARITY = 1'b1;
    defparam \CPU/PC[13]~FF .SR_SYNC = 1'b1;
    defparam \CPU/PC[13]~FF .SR_VALUE = 1'b0;
    defparam \CPU/PC[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/PC[14]~FF  (.D(\CPU/n2050 ), .CE(\CPU/state[2] ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\CPU/PC[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/PC[14]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/PC[14]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/PC[14]~FF .SR_POLARITY = 1'b0;
    defparam \CPU/PC[14]~FF .D_POLARITY = 1'b1;
    defparam \CPU/PC[14]~FF .SR_SYNC = 1'b1;
    defparam \CPU/PC[14]~FF .SR_VALUE = 1'b0;
    defparam \CPU/PC[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/PC[15]~FF  (.D(\CPU/n2049 ), .CE(\CPU/state[2] ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\CPU/PC[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/PC[15]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/PC[15]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/PC[15]~FF .SR_POLARITY = 1'b0;
    defparam \CPU/PC[15]~FF .D_POLARITY = 1'b1;
    defparam \CPU/PC[15]~FF .SR_SYNC = 1'b1;
    defparam \CPU/PC[15]~FF .SR_VALUE = 1'b0;
    defparam \CPU/PC[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/PC[16]~FF  (.D(\CPU/n2048 ), .CE(\CPU/state[2] ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\CPU/PC[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/PC[16]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/PC[16]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/PC[16]~FF .SR_POLARITY = 1'b0;
    defparam \CPU/PC[16]~FF .D_POLARITY = 1'b1;
    defparam \CPU/PC[16]~FF .SR_SYNC = 1'b1;
    defparam \CPU/PC[16]~FF .SR_VALUE = 1'b0;
    defparam \CPU/PC[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/PC[17]~FF  (.D(\CPU/n2047 ), .CE(\CPU/state[2] ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\CPU/PC[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/PC[17]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/PC[17]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/PC[17]~FF .SR_POLARITY = 1'b0;
    defparam \CPU/PC[17]~FF .D_POLARITY = 1'b1;
    defparam \CPU/PC[17]~FF .SR_SYNC = 1'b1;
    defparam \CPU/PC[17]~FF .SR_VALUE = 1'b0;
    defparam \CPU/PC[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/PC[18]~FF  (.D(\CPU/n2046 ), .CE(\CPU/state[2] ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\CPU/PC[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/PC[18]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/PC[18]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/PC[18]~FF .SR_POLARITY = 1'b0;
    defparam \CPU/PC[18]~FF .D_POLARITY = 1'b1;
    defparam \CPU/PC[18]~FF .SR_SYNC = 1'b1;
    defparam \CPU/PC[18]~FF .SR_VALUE = 1'b0;
    defparam \CPU/PC[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/PC[19]~FF  (.D(\CPU/n2045 ), .CE(\CPU/state[2] ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\CPU/PC[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/PC[19]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/PC[19]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/PC[19]~FF .SR_POLARITY = 1'b0;
    defparam \CPU/PC[19]~FF .D_POLARITY = 1'b1;
    defparam \CPU/PC[19]~FF .SR_SYNC = 1'b1;
    defparam \CPU/PC[19]~FF .SR_VALUE = 1'b0;
    defparam \CPU/PC[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/PC[20]~FF  (.D(\CPU/n2044 ), .CE(\CPU/state[2] ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\CPU/PC[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/PC[20]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/PC[20]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/PC[20]~FF .SR_POLARITY = 1'b0;
    defparam \CPU/PC[20]~FF .D_POLARITY = 1'b1;
    defparam \CPU/PC[20]~FF .SR_SYNC = 1'b1;
    defparam \CPU/PC[20]~FF .SR_VALUE = 1'b0;
    defparam \CPU/PC[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/PC[21]~FF  (.D(\CPU/n2043 ), .CE(\CPU/state[2] ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\CPU/PC[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/PC[21]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/PC[21]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/PC[21]~FF .SR_POLARITY = 1'b0;
    defparam \CPU/PC[21]~FF .D_POLARITY = 1'b1;
    defparam \CPU/PC[21]~FF .SR_SYNC = 1'b1;
    defparam \CPU/PC[21]~FF .SR_VALUE = 1'b0;
    defparam \CPU/PC[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/PC[22]~FF  (.D(\CPU/n2042 ), .CE(\CPU/state[2] ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\CPU/PC[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/PC[22]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/PC[22]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/PC[22]~FF .SR_POLARITY = 1'b0;
    defparam \CPU/PC[22]~FF .D_POLARITY = 1'b1;
    defparam \CPU/PC[22]~FF .SR_SYNC = 1'b1;
    defparam \CPU/PC[22]~FF .SR_VALUE = 1'b0;
    defparam \CPU/PC[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/PC[23]~FF  (.D(\CPU/n2041 ), .CE(\CPU/state[2] ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\CPU/PC[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/PC[23]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/PC[23]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/PC[23]~FF .SR_POLARITY = 1'b0;
    defparam \CPU/PC[23]~FF .D_POLARITY = 1'b1;
    defparam \CPU/PC[23]~FF .SR_SYNC = 1'b1;
    defparam \CPU/PC[23]~FF .SR_VALUE = 1'b0;
    defparam \CPU/PC[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/instr[3]~FF  (.D(\mem_rdata[3] ), .CE(\CPU/n3447 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/instr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/instr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/instr[3]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/instr[3]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/instr[3]~FF .D_POLARITY = 1'b1;
    defparam \CPU/instr[3]~FF .SR_SYNC = 1'b1;
    defparam \CPU/instr[3]~FF .SR_VALUE = 1'b0;
    defparam \CPU/instr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/instr[4]~FF  (.D(\mem_rdata[4] ), .CE(\CPU/n3447 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/instr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/instr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/instr[4]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/instr[4]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/instr[4]~FF .D_POLARITY = 1'b1;
    defparam \CPU/instr[4]~FF .SR_SYNC = 1'b1;
    defparam \CPU/instr[4]~FF .SR_VALUE = 1'b0;
    defparam \CPU/instr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/instr[5]~FF  (.D(\mem_rdata[5] ), .CE(\CPU/n3447 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/instr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/instr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/instr[5]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/instr[5]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/instr[5]~FF .D_POLARITY = 1'b1;
    defparam \CPU/instr[5]~FF .SR_SYNC = 1'b1;
    defparam \CPU/instr[5]~FF .SR_VALUE = 1'b0;
    defparam \CPU/instr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/instr[6]~FF  (.D(\mem_rdata[6] ), .CE(\CPU/n3447 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/instr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/instr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/instr[6]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/instr[6]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/instr[6]~FF .D_POLARITY = 1'b1;
    defparam \CPU/instr[6]~FF .SR_SYNC = 1'b1;
    defparam \CPU/instr[6]~FF .SR_VALUE = 1'b0;
    defparam \CPU/instr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/instr[7]~FF  (.D(\mem_rdata[7] ), .CE(\CPU/n3447 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/instr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/instr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/instr[7]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/instr[7]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/instr[7]~FF .D_POLARITY = 1'b1;
    defparam \CPU/instr[7]~FF .SR_SYNC = 1'b1;
    defparam \CPU/instr[7]~FF .SR_VALUE = 1'b0;
    defparam \CPU/instr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/instr[8]~FF  (.D(\mem_rdata[8] ), .CE(\CPU/n3447 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/instr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/instr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/instr[8]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/instr[8]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/instr[8]~FF .D_POLARITY = 1'b1;
    defparam \CPU/instr[8]~FF .SR_SYNC = 1'b1;
    defparam \CPU/instr[8]~FF .SR_VALUE = 1'b0;
    defparam \CPU/instr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/instr[9]~FF  (.D(\mem_rdata[9] ), .CE(\CPU/n3447 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/instr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/instr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/instr[9]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/instr[9]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/instr[9]~FF .D_POLARITY = 1'b1;
    defparam \CPU/instr[9]~FF .SR_SYNC = 1'b1;
    defparam \CPU/instr[9]~FF .SR_VALUE = 1'b0;
    defparam \CPU/instr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/instr[10]~FF  (.D(\mem_rdata[10] ), .CE(\CPU/n3447 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/instr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/instr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/instr[10]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/instr[10]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/instr[10]~FF .D_POLARITY = 1'b1;
    defparam \CPU/instr[10]~FF .SR_SYNC = 1'b1;
    defparam \CPU/instr[10]~FF .SR_VALUE = 1'b0;
    defparam \CPU/instr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/instr[11]~FF  (.D(\mem_rdata[11] ), .CE(\CPU/n3447 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/instr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/instr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/instr[11]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/instr[11]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/instr[11]~FF .D_POLARITY = 1'b1;
    defparam \CPU/instr[11]~FF .SR_SYNC = 1'b1;
    defparam \CPU/instr[11]~FF .SR_VALUE = 1'b0;
    defparam \CPU/instr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/instr[12]~FF  (.D(\mem_rdata[12] ), .CE(\CPU/n3447 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/instr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/instr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/instr[12]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/instr[12]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/instr[12]~FF .D_POLARITY = 1'b1;
    defparam \CPU/instr[12]~FF .SR_SYNC = 1'b1;
    defparam \CPU/instr[12]~FF .SR_VALUE = 1'b0;
    defparam \CPU/instr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/instr[13]~FF  (.D(\mem_rdata[13] ), .CE(\CPU/n3447 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/instr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/instr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/instr[13]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/instr[13]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/instr[13]~FF .D_POLARITY = 1'b1;
    defparam \CPU/instr[13]~FF .SR_SYNC = 1'b1;
    defparam \CPU/instr[13]~FF .SR_VALUE = 1'b0;
    defparam \CPU/instr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/instr[14]~FF  (.D(\mem_rdata[14] ), .CE(\CPU/n3447 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/instr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/instr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/instr[14]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/instr[14]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/instr[14]~FF .D_POLARITY = 1'b1;
    defparam \CPU/instr[14]~FF .SR_SYNC = 1'b1;
    defparam \CPU/instr[14]~FF .SR_VALUE = 1'b0;
    defparam \CPU/instr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/instr[15]~FF  (.D(\mem_rdata[15] ), .CE(\CPU/n3447 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/instr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/instr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/instr[15]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/instr[15]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/instr[15]~FF .D_POLARITY = 1'b1;
    defparam \CPU/instr[15]~FF .SR_SYNC = 1'b1;
    defparam \CPU/instr[15]~FF .SR_VALUE = 1'b0;
    defparam \CPU/instr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/instr[16]~FF  (.D(\mem_rdata[16] ), .CE(\CPU/n3447 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/instr[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/instr[16]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/instr[16]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/instr[16]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/instr[16]~FF .D_POLARITY = 1'b1;
    defparam \CPU/instr[16]~FF .SR_SYNC = 1'b1;
    defparam \CPU/instr[16]~FF .SR_VALUE = 1'b0;
    defparam \CPU/instr[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/instr[17]~FF  (.D(\mem_rdata[17] ), .CE(\CPU/n3447 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/instr[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/instr[17]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/instr[17]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/instr[17]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/instr[17]~FF .D_POLARITY = 1'b1;
    defparam \CPU/instr[17]~FF .SR_SYNC = 1'b1;
    defparam \CPU/instr[17]~FF .SR_VALUE = 1'b0;
    defparam \CPU/instr[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/instr[18]~FF  (.D(\mem_rdata[18] ), .CE(\CPU/n3447 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/instr[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/instr[18]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/instr[18]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/instr[18]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/instr[18]~FF .D_POLARITY = 1'b1;
    defparam \CPU/instr[18]~FF .SR_SYNC = 1'b1;
    defparam \CPU/instr[18]~FF .SR_VALUE = 1'b0;
    defparam \CPU/instr[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/instr[19]~FF  (.D(\mem_rdata[19] ), .CE(\CPU/n3447 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/instr[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/instr[19]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/instr[19]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/instr[19]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/instr[19]~FF .D_POLARITY = 1'b1;
    defparam \CPU/instr[19]~FF .SR_SYNC = 1'b1;
    defparam \CPU/instr[19]~FF .SR_VALUE = 1'b0;
    defparam \CPU/instr[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/instr[20]~FF  (.D(\mem_rdata[20] ), .CE(\CPU/n3447 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/instr[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/instr[20]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/instr[20]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/instr[20]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/instr[20]~FF .D_POLARITY = 1'b1;
    defparam \CPU/instr[20]~FF .SR_SYNC = 1'b1;
    defparam \CPU/instr[20]~FF .SR_VALUE = 1'b0;
    defparam \CPU/instr[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/instr[21]~FF  (.D(\mem_rdata[21] ), .CE(\CPU/n3447 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/instr[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/instr[21]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/instr[21]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/instr[21]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/instr[21]~FF .D_POLARITY = 1'b1;
    defparam \CPU/instr[21]~FF .SR_SYNC = 1'b1;
    defparam \CPU/instr[21]~FF .SR_VALUE = 1'b0;
    defparam \CPU/instr[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/instr[22]~FF  (.D(\mem_rdata[22] ), .CE(\CPU/n3447 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/instr[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/instr[22]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/instr[22]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/instr[22]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/instr[22]~FF .D_POLARITY = 1'b1;
    defparam \CPU/instr[22]~FF .SR_SYNC = 1'b1;
    defparam \CPU/instr[22]~FF .SR_VALUE = 1'b0;
    defparam \CPU/instr[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/instr[23]~FF  (.D(\mem_rdata[23] ), .CE(\CPU/n3447 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/instr[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/instr[23]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/instr[23]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/instr[23]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/instr[23]~FF .D_POLARITY = 1'b1;
    defparam \CPU/instr[23]~FF .SR_SYNC = 1'b1;
    defparam \CPU/instr[23]~FF .SR_VALUE = 1'b0;
    defparam \CPU/instr[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/instr[24]~FF  (.D(\mem_rdata[24] ), .CE(\CPU/n3447 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/instr[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/instr[24]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/instr[24]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/instr[24]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/instr[24]~FF .D_POLARITY = 1'b1;
    defparam \CPU/instr[24]~FF .SR_SYNC = 1'b1;
    defparam \CPU/instr[24]~FF .SR_VALUE = 1'b0;
    defparam \CPU/instr[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/instr[25]~FF  (.D(\mem_rdata[25] ), .CE(\CPU/n3447 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/instr[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/instr[25]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/instr[25]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/instr[25]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/instr[25]~FF .D_POLARITY = 1'b1;
    defparam \CPU/instr[25]~FF .SR_SYNC = 1'b1;
    defparam \CPU/instr[25]~FF .SR_VALUE = 1'b0;
    defparam \CPU/instr[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/instr[26]~FF  (.D(\mem_rdata[26] ), .CE(\CPU/n3447 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/instr[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/instr[26]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/instr[26]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/instr[26]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/instr[26]~FF .D_POLARITY = 1'b1;
    defparam \CPU/instr[26]~FF .SR_SYNC = 1'b1;
    defparam \CPU/instr[26]~FF .SR_VALUE = 1'b0;
    defparam \CPU/instr[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/instr[27]~FF  (.D(\mem_rdata[27] ), .CE(\CPU/n3447 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/instr[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/instr[27]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/instr[27]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/instr[27]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/instr[27]~FF .D_POLARITY = 1'b1;
    defparam \CPU/instr[27]~FF .SR_SYNC = 1'b1;
    defparam \CPU/instr[27]~FF .SR_VALUE = 1'b0;
    defparam \CPU/instr[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/instr[28]~FF  (.D(\mem_rdata[28] ), .CE(\CPU/n3447 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/instr[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/instr[28]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/instr[28]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/instr[28]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/instr[28]~FF .D_POLARITY = 1'b1;
    defparam \CPU/instr[28]~FF .SR_SYNC = 1'b1;
    defparam \CPU/instr[28]~FF .SR_VALUE = 1'b0;
    defparam \CPU/instr[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/instr[29]~FF  (.D(\mem_rdata[29] ), .CE(\CPU/n3447 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/instr[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/instr[29]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/instr[29]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/instr[29]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/instr[29]~FF .D_POLARITY = 1'b1;
    defparam \CPU/instr[29]~FF .SR_SYNC = 1'b1;
    defparam \CPU/instr[29]~FF .SR_VALUE = 1'b0;
    defparam \CPU/instr[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/instr[30]~FF  (.D(\mem_rdata[30] ), .CE(\CPU/n3447 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/instr[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/instr[30]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/instr[30]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/instr[30]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/instr[30]~FF .D_POLARITY = 1'b1;
    defparam \CPU/instr[30]~FF .SR_SYNC = 1'b1;
    defparam \CPU/instr[30]~FF .SR_VALUE = 1'b0;
    defparam \CPU/instr[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/instr[31]~FF  (.D(\mem_rdata[31] ), .CE(\CPU/n3447 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/instr[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/instr[31]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/instr[31]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/instr[31]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/instr[31]~FF .D_POLARITY = 1'b1;
    defparam \CPU/instr[31]~FF .SR_SYNC = 1'b1;
    defparam \CPU/instr[31]~FF .SR_VALUE = 1'b0;
    defparam \CPU/instr[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/cycles[1]~FF  (.D(n14), .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\CPU/cycles[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/cycles[1]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/cycles[1]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/cycles[1]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/cycles[1]~FF .D_POLARITY = 1'b1;
    defparam \CPU/cycles[1]~FF .SR_SYNC = 1'b1;
    defparam \CPU/cycles[1]~FF .SR_VALUE = 1'b0;
    defparam \CPU/cycles[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/cycles[2]~FF  (.D(n567), .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\CPU/cycles[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/cycles[2]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/cycles[2]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/cycles[2]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/cycles[2]~FF .D_POLARITY = 1'b1;
    defparam \CPU/cycles[2]~FF .SR_SYNC = 1'b1;
    defparam \CPU/cycles[2]~FF .SR_VALUE = 1'b0;
    defparam \CPU/cycles[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/cycles[3]~FF  (.D(n565), .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\CPU/cycles[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/cycles[3]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/cycles[3]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/cycles[3]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/cycles[3]~FF .D_POLARITY = 1'b1;
    defparam \CPU/cycles[3]~FF .SR_SYNC = 1'b1;
    defparam \CPU/cycles[3]~FF .SR_VALUE = 1'b0;
    defparam \CPU/cycles[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/cycles[4]~FF  (.D(n563), .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\CPU/cycles[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/cycles[4]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/cycles[4]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/cycles[4]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/cycles[4]~FF .D_POLARITY = 1'b1;
    defparam \CPU/cycles[4]~FF .SR_SYNC = 1'b1;
    defparam \CPU/cycles[4]~FF .SR_VALUE = 1'b0;
    defparam \CPU/cycles[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/cycles[5]~FF  (.D(n561), .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\CPU/cycles[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/cycles[5]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/cycles[5]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/cycles[5]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/cycles[5]~FF .D_POLARITY = 1'b1;
    defparam \CPU/cycles[5]~FF .SR_SYNC = 1'b1;
    defparam \CPU/cycles[5]~FF .SR_VALUE = 1'b0;
    defparam \CPU/cycles[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/cycles[6]~FF  (.D(n559), .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\CPU/cycles[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/cycles[6]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/cycles[6]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/cycles[6]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/cycles[6]~FF .D_POLARITY = 1'b1;
    defparam \CPU/cycles[6]~FF .SR_SYNC = 1'b1;
    defparam \CPU/cycles[6]~FF .SR_VALUE = 1'b0;
    defparam \CPU/cycles[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/cycles[7]~FF  (.D(n557), .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\CPU/cycles[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/cycles[7]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/cycles[7]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/cycles[7]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/cycles[7]~FF .D_POLARITY = 1'b1;
    defparam \CPU/cycles[7]~FF .SR_SYNC = 1'b1;
    defparam \CPU/cycles[7]~FF .SR_VALUE = 1'b0;
    defparam \CPU/cycles[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/cycles[8]~FF  (.D(n555), .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\CPU/cycles[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/cycles[8]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/cycles[8]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/cycles[8]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/cycles[8]~FF .D_POLARITY = 1'b1;
    defparam \CPU/cycles[8]~FF .SR_SYNC = 1'b1;
    defparam \CPU/cycles[8]~FF .SR_VALUE = 1'b0;
    defparam \CPU/cycles[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/cycles[9]~FF  (.D(n553), .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\CPU/cycles[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/cycles[9]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/cycles[9]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/cycles[9]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/cycles[9]~FF .D_POLARITY = 1'b1;
    defparam \CPU/cycles[9]~FF .SR_SYNC = 1'b1;
    defparam \CPU/cycles[9]~FF .SR_VALUE = 1'b0;
    defparam \CPU/cycles[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/cycles[10]~FF  (.D(n551), .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\CPU/cycles[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/cycles[10]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/cycles[10]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/cycles[10]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/cycles[10]~FF .D_POLARITY = 1'b1;
    defparam \CPU/cycles[10]~FF .SR_SYNC = 1'b1;
    defparam \CPU/cycles[10]~FF .SR_VALUE = 1'b0;
    defparam \CPU/cycles[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/cycles[11]~FF  (.D(n549), .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\CPU/cycles[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/cycles[11]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/cycles[11]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/cycles[11]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/cycles[11]~FF .D_POLARITY = 1'b1;
    defparam \CPU/cycles[11]~FF .SR_SYNC = 1'b1;
    defparam \CPU/cycles[11]~FF .SR_VALUE = 1'b0;
    defparam \CPU/cycles[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/cycles[12]~FF  (.D(n547), .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\CPU/cycles[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/cycles[12]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/cycles[12]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/cycles[12]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/cycles[12]~FF .D_POLARITY = 1'b1;
    defparam \CPU/cycles[12]~FF .SR_SYNC = 1'b1;
    defparam \CPU/cycles[12]~FF .SR_VALUE = 1'b0;
    defparam \CPU/cycles[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/cycles[13]~FF  (.D(n545), .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\CPU/cycles[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/cycles[13]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/cycles[13]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/cycles[13]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/cycles[13]~FF .D_POLARITY = 1'b1;
    defparam \CPU/cycles[13]~FF .SR_SYNC = 1'b1;
    defparam \CPU/cycles[13]~FF .SR_VALUE = 1'b0;
    defparam \CPU/cycles[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/cycles[14]~FF  (.D(n543), .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\CPU/cycles[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/cycles[14]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/cycles[14]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/cycles[14]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/cycles[14]~FF .D_POLARITY = 1'b1;
    defparam \CPU/cycles[14]~FF .SR_SYNC = 1'b1;
    defparam \CPU/cycles[14]~FF .SR_VALUE = 1'b0;
    defparam \CPU/cycles[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/cycles[15]~FF  (.D(n541), .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\CPU/cycles[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/cycles[15]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/cycles[15]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/cycles[15]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/cycles[15]~FF .D_POLARITY = 1'b1;
    defparam \CPU/cycles[15]~FF .SR_SYNC = 1'b1;
    defparam \CPU/cycles[15]~FF .SR_VALUE = 1'b0;
    defparam \CPU/cycles[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/cycles[16]~FF  (.D(n539), .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\CPU/cycles[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/cycles[16]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/cycles[16]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/cycles[16]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/cycles[16]~FF .D_POLARITY = 1'b1;
    defparam \CPU/cycles[16]~FF .SR_SYNC = 1'b1;
    defparam \CPU/cycles[16]~FF .SR_VALUE = 1'b0;
    defparam \CPU/cycles[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/cycles[17]~FF  (.D(n537), .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\CPU/cycles[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/cycles[17]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/cycles[17]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/cycles[17]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/cycles[17]~FF .D_POLARITY = 1'b1;
    defparam \CPU/cycles[17]~FF .SR_SYNC = 1'b1;
    defparam \CPU/cycles[17]~FF .SR_VALUE = 1'b0;
    defparam \CPU/cycles[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/cycles[18]~FF  (.D(n535), .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\CPU/cycles[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/cycles[18]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/cycles[18]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/cycles[18]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/cycles[18]~FF .D_POLARITY = 1'b1;
    defparam \CPU/cycles[18]~FF .SR_SYNC = 1'b1;
    defparam \CPU/cycles[18]~FF .SR_VALUE = 1'b0;
    defparam \CPU/cycles[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/cycles[19]~FF  (.D(n533), .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\CPU/cycles[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/cycles[19]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/cycles[19]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/cycles[19]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/cycles[19]~FF .D_POLARITY = 1'b1;
    defparam \CPU/cycles[19]~FF .SR_SYNC = 1'b1;
    defparam \CPU/cycles[19]~FF .SR_VALUE = 1'b0;
    defparam \CPU/cycles[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/cycles[20]~FF  (.D(n531), .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\CPU/cycles[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/cycles[20]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/cycles[20]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/cycles[20]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/cycles[20]~FF .D_POLARITY = 1'b1;
    defparam \CPU/cycles[20]~FF .SR_SYNC = 1'b1;
    defparam \CPU/cycles[20]~FF .SR_VALUE = 1'b0;
    defparam \CPU/cycles[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/cycles[21]~FF  (.D(n529), .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\CPU/cycles[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/cycles[21]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/cycles[21]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/cycles[21]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/cycles[21]~FF .D_POLARITY = 1'b1;
    defparam \CPU/cycles[21]~FF .SR_SYNC = 1'b1;
    defparam \CPU/cycles[21]~FF .SR_VALUE = 1'b0;
    defparam \CPU/cycles[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/cycles[22]~FF  (.D(n527), .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\CPU/cycles[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/cycles[22]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/cycles[22]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/cycles[22]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/cycles[22]~FF .D_POLARITY = 1'b1;
    defparam \CPU/cycles[22]~FF .SR_SYNC = 1'b1;
    defparam \CPU/cycles[22]~FF .SR_VALUE = 1'b0;
    defparam \CPU/cycles[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/cycles[23]~FF  (.D(n525), .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\CPU/cycles[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/cycles[23]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/cycles[23]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/cycles[23]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/cycles[23]~FF .D_POLARITY = 1'b1;
    defparam \CPU/cycles[23]~FF .SR_SYNC = 1'b1;
    defparam \CPU/cycles[23]~FF .SR_VALUE = 1'b0;
    defparam \CPU/cycles[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/cycles[24]~FF  (.D(n523), .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\CPU/cycles[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/cycles[24]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/cycles[24]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/cycles[24]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/cycles[24]~FF .D_POLARITY = 1'b1;
    defparam \CPU/cycles[24]~FF .SR_SYNC = 1'b1;
    defparam \CPU/cycles[24]~FF .SR_VALUE = 1'b0;
    defparam \CPU/cycles[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/cycles[25]~FF  (.D(n521), .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\CPU/cycles[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/cycles[25]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/cycles[25]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/cycles[25]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/cycles[25]~FF .D_POLARITY = 1'b1;
    defparam \CPU/cycles[25]~FF .SR_SYNC = 1'b1;
    defparam \CPU/cycles[25]~FF .SR_VALUE = 1'b0;
    defparam \CPU/cycles[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/cycles[26]~FF  (.D(n519), .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\CPU/cycles[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/cycles[26]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/cycles[26]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/cycles[26]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/cycles[26]~FF .D_POLARITY = 1'b1;
    defparam \CPU/cycles[26]~FF .SR_SYNC = 1'b1;
    defparam \CPU/cycles[26]~FF .SR_VALUE = 1'b0;
    defparam \CPU/cycles[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/cycles[27]~FF  (.D(n517), .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\CPU/cycles[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/cycles[27]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/cycles[27]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/cycles[27]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/cycles[27]~FF .D_POLARITY = 1'b1;
    defparam \CPU/cycles[27]~FF .SR_SYNC = 1'b1;
    defparam \CPU/cycles[27]~FF .SR_VALUE = 1'b0;
    defparam \CPU/cycles[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/cycles[28]~FF  (.D(n515), .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\CPU/cycles[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/cycles[28]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/cycles[28]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/cycles[28]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/cycles[28]~FF .D_POLARITY = 1'b1;
    defparam \CPU/cycles[28]~FF .SR_SYNC = 1'b1;
    defparam \CPU/cycles[28]~FF .SR_VALUE = 1'b0;
    defparam \CPU/cycles[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/cycles[29]~FF  (.D(n513), .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\CPU/cycles[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/cycles[29]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/cycles[29]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/cycles[29]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/cycles[29]~FF .D_POLARITY = 1'b1;
    defparam \CPU/cycles[29]~FF .SR_SYNC = 1'b1;
    defparam \CPU/cycles[29]~FF .SR_VALUE = 1'b0;
    defparam \CPU/cycles[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/cycles[30]~FF  (.D(n511), .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\CPU/cycles[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/cycles[30]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/cycles[30]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/cycles[30]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/cycles[30]~FF .D_POLARITY = 1'b1;
    defparam \CPU/cycles[30]~FF .SR_SYNC = 1'b1;
    defparam \CPU/cycles[30]~FF .SR_VALUE = 1'b0;
    defparam \CPU/cycles[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/cycles[31]~FF  (.D(n510), .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\CPU/cycles[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/cycles[31]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/cycles[31]~FF .CE_POLARITY = 1'b1;
    defparam \CPU/cycles[31]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/cycles[31]~FF .D_POLARITY = 1'b1;
    defparam \CPU/cycles[31]~FF .SR_SYNC = 1'b1;
    defparam \CPU/cycles[31]~FF .SR_VALUE = 1'b0;
    defparam \CPU/cycles[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/aluReg[2]~FF  (.D(\CPU/n1065 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluReg[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluReg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluReg[2]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluReg[2]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluReg[2]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluReg[2]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluReg[2]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluReg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/aluReg[3]~FF  (.D(\CPU/n1064 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluReg[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluReg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluReg[3]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluReg[3]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluReg[3]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluReg[3]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluReg[3]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluReg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/aluReg[4]~FF  (.D(\CPU/n1063 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluReg[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluReg[4]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluReg[4]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluReg[4]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluReg[4]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluReg[4]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluReg[4]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluReg[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/aluReg[5]~FF  (.D(\CPU/n1062 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluReg[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluReg[5]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluReg[5]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluReg[5]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluReg[5]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluReg[5]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluReg[5]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluReg[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/aluReg[6]~FF  (.D(\CPU/n1061 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluReg[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluReg[6]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluReg[6]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluReg[6]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluReg[6]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluReg[6]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluReg[6]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluReg[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/aluReg[7]~FF  (.D(\CPU/n1060 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluReg[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluReg[7]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluReg[7]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluReg[7]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluReg[7]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluReg[7]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluReg[7]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluReg[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/aluReg[8]~FF  (.D(\CPU/n1059 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluReg[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluReg[8]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluReg[8]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluReg[8]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluReg[8]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluReg[8]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluReg[8]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluReg[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/aluReg[9]~FF  (.D(\CPU/n1058 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluReg[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluReg[9]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluReg[9]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluReg[9]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluReg[9]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluReg[9]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluReg[9]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluReg[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/aluReg[10]~FF  (.D(\CPU/n1057 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluReg[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluReg[10]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluReg[10]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluReg[10]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluReg[10]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluReg[10]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluReg[10]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluReg[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/aluReg[11]~FF  (.D(\CPU/n1056 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluReg[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluReg[11]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluReg[11]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluReg[11]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluReg[11]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluReg[11]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluReg[11]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluReg[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/aluReg[12]~FF  (.D(\CPU/n1055 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluReg[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluReg[12]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluReg[12]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluReg[12]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluReg[12]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluReg[12]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluReg[12]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluReg[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/aluReg[13]~FF  (.D(\CPU/n1054 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluReg[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluReg[13]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluReg[13]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluReg[13]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluReg[13]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluReg[13]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluReg[13]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluReg[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/aluReg[14]~FF  (.D(\CPU/n1053 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluReg[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluReg[14]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluReg[14]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluReg[14]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluReg[14]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluReg[14]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluReg[14]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluReg[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/aluReg[15]~FF  (.D(\CPU/n1052 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluReg[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluReg[15]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluReg[15]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluReg[15]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluReg[15]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluReg[15]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluReg[15]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluReg[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/aluReg[16]~FF  (.D(\CPU/n1051 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluReg[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluReg[16]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluReg[16]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluReg[16]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluReg[16]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluReg[16]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluReg[16]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluReg[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/aluReg[17]~FF  (.D(\CPU/n1050 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluReg[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluReg[17]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluReg[17]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluReg[17]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluReg[17]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluReg[17]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluReg[17]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluReg[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/aluReg[18]~FF  (.D(\CPU/n1049 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluReg[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluReg[18]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluReg[18]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluReg[18]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluReg[18]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluReg[18]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluReg[18]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluReg[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/aluReg[19]~FF  (.D(\CPU/n1048 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluReg[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluReg[19]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluReg[19]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluReg[19]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluReg[19]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluReg[19]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluReg[19]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluReg[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/aluReg[20]~FF  (.D(\CPU/n1047 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluReg[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluReg[20]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluReg[20]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluReg[20]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluReg[20]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluReg[20]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluReg[20]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluReg[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/aluReg[21]~FF  (.D(\CPU/n1046 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluReg[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluReg[21]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluReg[21]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluReg[21]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluReg[21]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluReg[21]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluReg[21]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluReg[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/aluReg[22]~FF  (.D(\CPU/n1045 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluReg[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluReg[22]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluReg[22]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluReg[22]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluReg[22]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluReg[22]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluReg[22]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluReg[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/aluReg[23]~FF  (.D(\CPU/n1044 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluReg[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluReg[23]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluReg[23]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluReg[23]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluReg[23]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluReg[23]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluReg[23]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluReg[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/aluReg[24]~FF  (.D(\CPU/n1043 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluReg[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluReg[24]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluReg[24]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluReg[24]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluReg[24]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluReg[24]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluReg[24]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluReg[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/aluReg[25]~FF  (.D(\CPU/n1042 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluReg[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluReg[25]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluReg[25]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluReg[25]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluReg[25]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluReg[25]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluReg[25]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluReg[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/aluReg[26]~FF  (.D(\CPU/n1041 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluReg[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluReg[26]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluReg[26]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluReg[26]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluReg[26]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluReg[26]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluReg[26]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluReg[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/aluReg[27]~FF  (.D(\CPU/n1040 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluReg[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluReg[27]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluReg[27]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluReg[27]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluReg[27]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluReg[27]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluReg[27]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluReg[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/aluReg[28]~FF  (.D(\CPU/n1039 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluReg[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluReg[28]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluReg[28]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluReg[28]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluReg[28]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluReg[28]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluReg[28]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluReg[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/aluReg[29]~FF  (.D(\CPU/n1038 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluReg[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluReg[29]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluReg[29]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluReg[29]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluReg[29]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluReg[29]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluReg[29]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluReg[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/aluReg[30]~FF  (.D(\CPU/n1037 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluReg[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluReg[30]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluReg[30]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluReg[30]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluReg[30]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluReg[30]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluReg[30]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluReg[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/aluReg[31]~FF  (.D(\CPU/n1036 ), .CE(ceg_net77), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/aluReg[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(178)
    defparam \CPU/aluReg[31]~FF .CLK_POLARITY = 1'b1;
    defparam \CPU/aluReg[31]~FF .CE_POLARITY = 1'b0;
    defparam \CPU/aluReg[31]~FF .SR_POLARITY = 1'b1;
    defparam \CPU/aluReg[31]~FF .D_POLARITY = 1'b1;
    defparam \CPU/aluReg[31]~FF .SR_SYNC = 1'b1;
    defparam \CPU/aluReg[31]~FF .SR_VALUE = 1'b0;
    defparam \CPU/aluReg[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart_ctrl[0]~FF  (.D(\mem_wdata[0] ), .CE(\per_uart/n25 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/uart_ctrl[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/perip_uart.v(42)
    defparam \per_uart/uart_ctrl[0]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart_ctrl[0]~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/uart_ctrl[0]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/uart_ctrl[0]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart_ctrl[0]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart_ctrl[0]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart_ctrl[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_dout[0]~FF  (.D(\per_uart/select_21/Select_0/n3 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_dout[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/perip_uart.v(51)
    defparam \uart_dout[0]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_dout[0]~FF .CE_POLARITY = 1'b1;
    defparam \uart_dout[0]~FF .SR_POLARITY = 1'b1;
    defparam \uart_dout[0]~FF .D_POLARITY = 1'b1;
    defparam \uart_dout[0]~FF .SR_SYNC = 1'b1;
    defparam \uart_dout[0]~FF .SR_VALUE = 1'b0;
    defparam \uart_dout[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/d_in_uart[0]~FF  (.D(\mem_wdata[0] ), .CE(\per_uart/n15 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/d_in_uart[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/perip_uart.v(42)
    defparam \per_uart/d_in_uart[0]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/d_in_uart[0]~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/d_in_uart[0]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/d_in_uart[0]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/d_in_uart[0]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/d_in_uart[0]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/d_in_uart[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart_ctrl[1]~FF  (.D(\mem_wdata[1] ), .CE(\per_uart/n25 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/uart_ctrl[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/perip_uart.v(42)
    defparam \per_uart/uart_ctrl[1]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart_ctrl[1]~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/uart_ctrl[1]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/uart_ctrl[1]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart_ctrl[1]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart_ctrl[1]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart_ctrl[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \LEDS~FF  (.D(\mem_wdata[2] ), .CE(\per_uart/n25 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(LEDS)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/perip_uart.v(42)
    defparam \LEDS~FF .CLK_POLARITY = 1'b1;
    defparam \LEDS~FF .CE_POLARITY = 1'b1;
    defparam \LEDS~FF .SR_POLARITY = 1'b1;
    defparam \LEDS~FF .D_POLARITY = 1'b1;
    defparam \LEDS~FF .SR_SYNC = 1'b1;
    defparam \LEDS~FF .SR_VALUE = 1'b0;
    defparam \LEDS~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_dout[1]~FF  (.D(\per_uart/select_21/Select_1/n3 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_dout[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/perip_uart.v(51)
    defparam \uart_dout[1]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_dout[1]~FF .CE_POLARITY = 1'b1;
    defparam \uart_dout[1]~FF .SR_POLARITY = 1'b1;
    defparam \uart_dout[1]~FF .D_POLARITY = 1'b1;
    defparam \uart_dout[1]~FF .SR_SYNC = 1'b1;
    defparam \uart_dout[1]~FF .SR_VALUE = 1'b0;
    defparam \uart_dout[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_dout[2]~FF  (.D(\per_uart/select_21/Select_2/n3 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_dout[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/perip_uart.v(51)
    defparam \uart_dout[2]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_dout[2]~FF .CE_POLARITY = 1'b1;
    defparam \uart_dout[2]~FF .SR_POLARITY = 1'b1;
    defparam \uart_dout[2]~FF .D_POLARITY = 1'b1;
    defparam \uart_dout[2]~FF .SR_SYNC = 1'b1;
    defparam \uart_dout[2]~FF .SR_VALUE = 1'b0;
    defparam \uart_dout[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_dout[3]~FF  (.D(\per_uart/select_21/Select_3/n3 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_dout[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/perip_uart.v(51)
    defparam \uart_dout[3]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_dout[3]~FF .CE_POLARITY = 1'b1;
    defparam \uart_dout[3]~FF .SR_POLARITY = 1'b1;
    defparam \uart_dout[3]~FF .D_POLARITY = 1'b1;
    defparam \uart_dout[3]~FF .SR_SYNC = 1'b1;
    defparam \uart_dout[3]~FF .SR_VALUE = 1'b0;
    defparam \uart_dout[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_dout[4]~FF  (.D(\per_uart/select_21/Select_4/n3 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_dout[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/perip_uart.v(51)
    defparam \uart_dout[4]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_dout[4]~FF .CE_POLARITY = 1'b1;
    defparam \uart_dout[4]~FF .SR_POLARITY = 1'b1;
    defparam \uart_dout[4]~FF .D_POLARITY = 1'b1;
    defparam \uart_dout[4]~FF .SR_SYNC = 1'b1;
    defparam \uart_dout[4]~FF .SR_VALUE = 1'b0;
    defparam \uart_dout[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_dout[5]~FF  (.D(\per_uart/select_21/Select_5/n3 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_dout[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/perip_uart.v(51)
    defparam \uart_dout[5]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_dout[5]~FF .CE_POLARITY = 1'b1;
    defparam \uart_dout[5]~FF .SR_POLARITY = 1'b1;
    defparam \uart_dout[5]~FF .D_POLARITY = 1'b1;
    defparam \uart_dout[5]~FF .SR_SYNC = 1'b1;
    defparam \uart_dout[5]~FF .SR_VALUE = 1'b0;
    defparam \uart_dout[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_dout[6]~FF  (.D(\per_uart/select_21/Select_6/n3 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_dout[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/perip_uart.v(51)
    defparam \uart_dout[6]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_dout[6]~FF .CE_POLARITY = 1'b1;
    defparam \uart_dout[6]~FF .SR_POLARITY = 1'b1;
    defparam \uart_dout[6]~FF .D_POLARITY = 1'b1;
    defparam \uart_dout[6]~FF .SR_SYNC = 1'b1;
    defparam \uart_dout[6]~FF .SR_VALUE = 1'b0;
    defparam \uart_dout[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_dout[7]~FF  (.D(\per_uart/select_21/Select_7/n4 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_dout[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/perip_uart.v(51)
    defparam \uart_dout[7]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_dout[7]~FF .CE_POLARITY = 1'b1;
    defparam \uart_dout[7]~FF .SR_POLARITY = 1'b1;
    defparam \uart_dout[7]~FF .D_POLARITY = 1'b1;
    defparam \uart_dout[7]~FF .SR_SYNC = 1'b1;
    defparam \uart_dout[7]~FF .SR_VALUE = 1'b0;
    defparam \uart_dout[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_dout[8]~FF  (.D(\per_uart/select_21/Select_8/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_dout[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/perip_uart.v(51)
    defparam \uart_dout[8]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_dout[8]~FF .CE_POLARITY = 1'b1;
    defparam \uart_dout[8]~FF .SR_POLARITY = 1'b1;
    defparam \uart_dout[8]~FF .D_POLARITY = 1'b1;
    defparam \uart_dout[8]~FF .SR_SYNC = 1'b1;
    defparam \uart_dout[8]~FF .SR_VALUE = 1'b0;
    defparam \uart_dout[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_dout[9]~FF  (.D(\per_uart/select_21/Select_9/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_dout[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/perip_uart.v(51)
    defparam \uart_dout[9]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_dout[9]~FF .CE_POLARITY = 1'b1;
    defparam \uart_dout[9]~FF .SR_POLARITY = 1'b1;
    defparam \uart_dout[9]~FF .D_POLARITY = 1'b1;
    defparam \uart_dout[9]~FF .SR_SYNC = 1'b1;
    defparam \uart_dout[9]~FF .SR_VALUE = 1'b0;
    defparam \uart_dout[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/uart_rxd1~FF  (.D(RXD), .CE(1'b1), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\per_uart/uart0/uart_rxd1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(56)
    defparam \per_uart/uart0/uart_rxd1~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/uart_rxd1~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/uart0/uart_rxd1~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/uart0/uart_rxd1~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/uart_rxd1~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/uart_rxd1~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/uart_rxd1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/uart_rxd2~FF  (.D(\per_uart/uart0/uart_rxd1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/uart0/uart_rxd2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(56)
    defparam \per_uart/uart0/uart_rxd2~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/uart_rxd2~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/uart0/uart_rxd2~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/uart0/uart_rxd2~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/uart_rxd2~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/uart_rxd2~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/uart_rxd2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/rx_busy~FF  (.D(\per_uart/uart0/n190 ), .CE(ceg_net530), 
           .CLK(\clk~O ), .SR(resetn), .Q(\per_uart/uart0/rx_busy )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(113)
    defparam \per_uart/uart0/rx_busy~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/rx_busy~FF .CE_POLARITY = 1'b0;
    defparam \per_uart/uart0/rx_busy~FF .SR_POLARITY = 1'b0;
    defparam \per_uart/uart0/rx_busy~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/rx_busy~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/rx_busy~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/rx_busy~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/rx_count16[0]~FF  (.D(\per_uart/uart0/n195 ), .CE(ceg_net176), 
           .CLK(\clk~O ), .SR(resetn), .Q(\per_uart/uart0/rx_count16[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(113)
    defparam \per_uart/uart0/rx_count16[0]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/rx_count16[0]~FF .CE_POLARITY = 1'b0;
    defparam \per_uart/uart0/rx_count16[0]~FF .SR_POLARITY = 1'b0;
    defparam \per_uart/uart0/rx_count16[0]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/rx_count16[0]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/rx_count16[0]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/rx_count16[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/rx_bitcount[0]~FF  (.D(\per_uart/uart0/n200 ), 
           .CE(ceg_net530), .CLK(\clk~O ), .SR(resetn), .Q(\per_uart/uart0/rx_bitcount[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(113)
    defparam \per_uart/uart0/rx_bitcount[0]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/rx_bitcount[0]~FF .CE_POLARITY = 1'b0;
    defparam \per_uart/uart0/rx_bitcount[0]~FF .SR_POLARITY = 1'b0;
    defparam \per_uart/uart0/rx_bitcount[0]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/rx_bitcount[0]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/rx_bitcount[0]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/rx_bitcount[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/rx_data[0]~FF  (.D(\per_uart/uart0/rxd_reg[0] ), .CE(\per_uart/uart0/n581 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/rx_data[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(113)
    defparam \per_uart/rx_data[0]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/rx_data[0]~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/rx_data[0]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/rx_data[0]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/rx_data[0]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/rx_data[0]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/rx_data[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/rx_avail~FF  (.D(\per_uart/uart0/n576 ), .CE(ceg_net140), 
           .CLK(\clk~O ), .SR(resetn), .Q(\per_uart/rx_avail )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(113)
    defparam \per_uart/rx_avail~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/rx_avail~FF .CE_POLARITY = 1'b0;
    defparam \per_uart/rx_avail~FF .SR_POLARITY = 1'b0;
    defparam \per_uart/rx_avail~FF .D_POLARITY = 1'b1;
    defparam \per_uart/rx_avail~FF .SR_SYNC = 1'b1;
    defparam \per_uart/rx_avail~FF .SR_VALUE = 1'b0;
    defparam \per_uart/rx_avail~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/rx_error~FF  (.D(\per_uart/uart0/n242 ), .CE(ceg_net144), 
           .CLK(\clk~O ), .SR(resetn), .Q(\per_uart/rx_error )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(113)
    defparam \per_uart/rx_error~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/rx_error~FF .CE_POLARITY = 1'b0;
    defparam \per_uart/rx_error~FF .SR_POLARITY = 1'b0;
    defparam \per_uart/rx_error~FF .D_POLARITY = 1'b1;
    defparam \per_uart/rx_error~FF .SR_SYNC = 1'b1;
    defparam \per_uart/rx_error~FF .SR_VALUE = 1'b0;
    defparam \per_uart/rx_error~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/rxd_reg[0]~FF  (.D(\per_uart/uart0/rxd_reg[1] ), 
           .CE(\per_uart/uart0/n582 ), .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/uart0/rxd_reg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(113)
    defparam \per_uart/uart0/rxd_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/rxd_reg[0]~FF .CE_POLARITY = 1'b0;
    defparam \per_uart/uart0/rxd_reg[0]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/uart0/rxd_reg[0]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/rxd_reg[0]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/rxd_reg[0]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/rxd_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/tx_busy~FF  (.D(1'b1), .CE(\per_uart/uart0/n316 ), 
           .CLK(\clk~O ), .SR(\per_uart/uart0/n601 ), .Q(\per_uart/tx_busy )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(157)
    defparam \per_uart/tx_busy~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/tx_busy~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/tx_busy~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/tx_busy~FF .D_POLARITY = 1'b1;
    defparam \per_uart/tx_busy~FF .SR_SYNC = 1'b1;
    defparam \per_uart/tx_busy~FF .SR_VALUE = 1'b0;
    defparam \per_uart/tx_busy~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/tx_count16[0]~FF  (.D(\per_uart/uart0/n422 ), .CE(ceg_net203), 
           .CLK(\clk~O ), .SR(resetn), .Q(\per_uart/uart0/tx_count16[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(157)
    defparam \per_uart/uart0/tx_count16[0]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/tx_count16[0]~FF .CE_POLARITY = 1'b0;
    defparam \per_uart/uart0/tx_count16[0]~FF .SR_POLARITY = 1'b0;
    defparam \per_uart/uart0/tx_count16[0]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/tx_count16[0]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/tx_count16[0]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/tx_count16[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \TXD~FF  (.D(\per_uart/uart0/n386 ), .CE(ceg_net155), .CLK(\clk~O ), 
           .SR(resetn), .Q(TXD)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(157)
    defparam \TXD~FF .CLK_POLARITY = 1'b1;
    defparam \TXD~FF .CE_POLARITY = 1'b1;
    defparam \TXD~FF .SR_POLARITY = 1'b0;
    defparam \TXD~FF .D_POLARITY = 1'b1;
    defparam \TXD~FF .SR_SYNC = 1'b1;
    defparam \TXD~FF .SR_VALUE = 1'b1;
    defparam \TXD~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/txd_reg[0]~FF  (.D(\per_uart/uart0/n438 ), .CE(ceg_net159), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/uart0/txd_reg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(157)
    defparam \per_uart/uart0/txd_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/txd_reg[0]~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/uart0/txd_reg[0]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/uart0/txd_reg[0]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/txd_reg[0]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/txd_reg[0]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/txd_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/tx_bitcount[0]~FF  (.D(\per_uart/uart0/n427 ), 
           .CE(ceg_net246), .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/uart0/tx_bitcount[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(157)
    defparam \per_uart/uart0/tx_bitcount[0]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/tx_bitcount[0]~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/uart0/tx_bitcount[0]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/uart0/tx_bitcount[0]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/tx_bitcount[0]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/tx_bitcount[0]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/tx_bitcount[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/enable16_counter[0]~FF  (.D(\per_uart/uart0/enable16_counter[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\per_uart/uart0/n552 ), .Q(\per_uart/uart0/enable16_counter[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(44)
    defparam \per_uart/uart0/enable16_counter[0]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/enable16_counter[0]~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/uart0/enable16_counter[0]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/uart0/enable16_counter[0]~FF .D_POLARITY = 1'b0;
    defparam \per_uart/uart0/enable16_counter[0]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/enable16_counter[0]~FF .SR_VALUE = 1'b1;
    defparam \per_uart/uart0/enable16_counter[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/rx_count16[1]~FF  (.D(\per_uart/uart0/n194 ), .CE(ceg_net176), 
           .CLK(\clk~O ), .SR(resetn), .Q(\per_uart/uart0/rx_count16[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(113)
    defparam \per_uart/uart0/rx_count16[1]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/rx_count16[1]~FF .CE_POLARITY = 1'b0;
    defparam \per_uart/uart0/rx_count16[1]~FF .SR_POLARITY = 1'b0;
    defparam \per_uart/uart0/rx_count16[1]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/rx_count16[1]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/rx_count16[1]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/rx_count16[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/rx_count16[2]~FF  (.D(\per_uart/uart0/n193 ), .CE(ceg_net176), 
           .CLK(\clk~O ), .SR(resetn), .Q(\per_uart/uart0/rx_count16[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(113)
    defparam \per_uart/uart0/rx_count16[2]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/rx_count16[2]~FF .CE_POLARITY = 1'b0;
    defparam \per_uart/uart0/rx_count16[2]~FF .SR_POLARITY = 1'b0;
    defparam \per_uart/uart0/rx_count16[2]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/rx_count16[2]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/rx_count16[2]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/rx_count16[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/rx_count16[3]~FF  (.D(\per_uart/uart0/n192 ), .CE(ceg_net176), 
           .CLK(\clk~O ), .SR(resetn), .Q(\per_uart/uart0/rx_count16[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(113)
    defparam \per_uart/uart0/rx_count16[3]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/rx_count16[3]~FF .CE_POLARITY = 1'b0;
    defparam \per_uart/uart0/rx_count16[3]~FF .SR_POLARITY = 1'b0;
    defparam \per_uart/uart0/rx_count16[3]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/rx_count16[3]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/rx_count16[3]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/rx_count16[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/rx_bitcount[1]~FF  (.D(\per_uart/uart0/n199 ), 
           .CE(ceg_net530), .CLK(\clk~O ), .SR(resetn), .Q(\per_uart/uart0/rx_bitcount[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(113)
    defparam \per_uart/uart0/rx_bitcount[1]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/rx_bitcount[1]~FF .CE_POLARITY = 1'b0;
    defparam \per_uart/uart0/rx_bitcount[1]~FF .SR_POLARITY = 1'b0;
    defparam \per_uart/uart0/rx_bitcount[1]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/rx_bitcount[1]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/rx_bitcount[1]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/rx_bitcount[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/rx_bitcount[2]~FF  (.D(\per_uart/uart0/n198 ), 
           .CE(ceg_net530), .CLK(\clk~O ), .SR(resetn), .Q(\per_uart/uart0/rx_bitcount[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(113)
    defparam \per_uart/uart0/rx_bitcount[2]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/rx_bitcount[2]~FF .CE_POLARITY = 1'b0;
    defparam \per_uart/uart0/rx_bitcount[2]~FF .SR_POLARITY = 1'b0;
    defparam \per_uart/uart0/rx_bitcount[2]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/rx_bitcount[2]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/rx_bitcount[2]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/rx_bitcount[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/rx_bitcount[3]~FF  (.D(\per_uart/uart0/n197 ), 
           .CE(ceg_net530), .CLK(\clk~O ), .SR(resetn), .Q(\per_uart/uart0/rx_bitcount[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(113)
    defparam \per_uart/uart0/rx_bitcount[3]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/rx_bitcount[3]~FF .CE_POLARITY = 1'b0;
    defparam \per_uart/uart0/rx_bitcount[3]~FF .SR_POLARITY = 1'b0;
    defparam \per_uart/uart0/rx_bitcount[3]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/rx_bitcount[3]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/rx_bitcount[3]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/rx_bitcount[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/rx_data[1]~FF  (.D(\per_uart/uart0/rxd_reg[1] ), .CE(\per_uart/uart0/n581 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/rx_data[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(113)
    defparam \per_uart/rx_data[1]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/rx_data[1]~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/rx_data[1]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/rx_data[1]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/rx_data[1]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/rx_data[1]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/rx_data[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/rx_data[2]~FF  (.D(\per_uart/uart0/rxd_reg[2] ), .CE(\per_uart/uart0/n581 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/rx_data[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(113)
    defparam \per_uart/rx_data[2]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/rx_data[2]~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/rx_data[2]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/rx_data[2]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/rx_data[2]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/rx_data[2]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/rx_data[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/rx_data[3]~FF  (.D(\per_uart/uart0/rxd_reg[3] ), .CE(\per_uart/uart0/n581 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/rx_data[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(113)
    defparam \per_uart/rx_data[3]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/rx_data[3]~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/rx_data[3]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/rx_data[3]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/rx_data[3]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/rx_data[3]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/rx_data[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/rx_data[4]~FF  (.D(\per_uart/uart0/rxd_reg[4] ), .CE(\per_uart/uart0/n581 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/rx_data[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(113)
    defparam \per_uart/rx_data[4]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/rx_data[4]~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/rx_data[4]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/rx_data[4]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/rx_data[4]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/rx_data[4]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/rx_data[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/rx_data[5]~FF  (.D(\per_uart/uart0/rxd_reg[5] ), .CE(\per_uart/uart0/n581 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/rx_data[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(113)
    defparam \per_uart/rx_data[5]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/rx_data[5]~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/rx_data[5]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/rx_data[5]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/rx_data[5]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/rx_data[5]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/rx_data[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/rx_data[6]~FF  (.D(\per_uart/uart0/rxd_reg[6] ), .CE(\per_uart/uart0/n581 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/rx_data[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(113)
    defparam \per_uart/rx_data[6]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/rx_data[6]~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/rx_data[6]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/rx_data[6]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/rx_data[6]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/rx_data[6]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/rx_data[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/rx_data[7]~FF  (.D(\per_uart/uart0/rxd_reg[7] ), .CE(\per_uart/uart0/n581 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/rx_data[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(113)
    defparam \per_uart/rx_data[7]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/rx_data[7]~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/rx_data[7]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/rx_data[7]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/rx_data[7]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/rx_data[7]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/rx_data[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/rxd_reg[1]~FF  (.D(\per_uart/uart0/rxd_reg[2] ), 
           .CE(\per_uart/uart0/n582 ), .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/uart0/rxd_reg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(113)
    defparam \per_uart/uart0/rxd_reg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/rxd_reg[1]~FF .CE_POLARITY = 1'b0;
    defparam \per_uart/uart0/rxd_reg[1]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/uart0/rxd_reg[1]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/rxd_reg[1]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/rxd_reg[1]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/rxd_reg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/rxd_reg[2]~FF  (.D(\per_uart/uart0/rxd_reg[3] ), 
           .CE(\per_uart/uart0/n582 ), .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/uart0/rxd_reg[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(113)
    defparam \per_uart/uart0/rxd_reg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/rxd_reg[2]~FF .CE_POLARITY = 1'b0;
    defparam \per_uart/uart0/rxd_reg[2]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/uart0/rxd_reg[2]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/rxd_reg[2]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/rxd_reg[2]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/rxd_reg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/rxd_reg[3]~FF  (.D(\per_uart/uart0/rxd_reg[4] ), 
           .CE(\per_uart/uart0/n582 ), .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/uart0/rxd_reg[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(113)
    defparam \per_uart/uart0/rxd_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/rxd_reg[3]~FF .CE_POLARITY = 1'b0;
    defparam \per_uart/uart0/rxd_reg[3]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/uart0/rxd_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/rxd_reg[3]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/rxd_reg[3]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/rxd_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/rxd_reg[4]~FF  (.D(\per_uart/uart0/rxd_reg[5] ), 
           .CE(\per_uart/uart0/n582 ), .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/uart0/rxd_reg[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(113)
    defparam \per_uart/uart0/rxd_reg[4]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/rxd_reg[4]~FF .CE_POLARITY = 1'b0;
    defparam \per_uart/uart0/rxd_reg[4]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/uart0/rxd_reg[4]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/rxd_reg[4]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/rxd_reg[4]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/rxd_reg[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/rxd_reg[5]~FF  (.D(\per_uart/uart0/rxd_reg[6] ), 
           .CE(\per_uart/uart0/n582 ), .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/uart0/rxd_reg[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(113)
    defparam \per_uart/uart0/rxd_reg[5]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/rxd_reg[5]~FF .CE_POLARITY = 1'b0;
    defparam \per_uart/uart0/rxd_reg[5]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/uart0/rxd_reg[5]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/rxd_reg[5]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/rxd_reg[5]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/rxd_reg[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/rxd_reg[6]~FF  (.D(\per_uart/uart0/rxd_reg[7] ), 
           .CE(\per_uart/uart0/n582 ), .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/uart0/rxd_reg[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(113)
    defparam \per_uart/uart0/rxd_reg[6]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/rxd_reg[6]~FF .CE_POLARITY = 1'b0;
    defparam \per_uart/uart0/rxd_reg[6]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/uart0/rxd_reg[6]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/rxd_reg[6]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/rxd_reg[6]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/rxd_reg[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/rxd_reg[7]~FF  (.D(\per_uart/uart0/uart_rxd2 ), 
           .CE(\per_uart/uart0/n582 ), .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/uart0/rxd_reg[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(113)
    defparam \per_uart/uart0/rxd_reg[7]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/rxd_reg[7]~FF .CE_POLARITY = 1'b0;
    defparam \per_uart/uart0/rxd_reg[7]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/uart0/rxd_reg[7]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/rxd_reg[7]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/rxd_reg[7]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/rxd_reg[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/tx_count16[1]~FF  (.D(\per_uart/uart0/n421 ), .CE(ceg_net203), 
           .CLK(\clk~O ), .SR(resetn), .Q(\per_uart/uart0/tx_count16[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(157)
    defparam \per_uart/uart0/tx_count16[1]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/tx_count16[1]~FF .CE_POLARITY = 1'b0;
    defparam \per_uart/uart0/tx_count16[1]~FF .SR_POLARITY = 1'b0;
    defparam \per_uart/uart0/tx_count16[1]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/tx_count16[1]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/tx_count16[1]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/tx_count16[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/tx_count16[2]~FF  (.D(\per_uart/uart0/n420 ), .CE(ceg_net203), 
           .CLK(\clk~O ), .SR(resetn), .Q(\per_uart/uart0/tx_count16[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(157)
    defparam \per_uart/uart0/tx_count16[2]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/tx_count16[2]~FF .CE_POLARITY = 1'b0;
    defparam \per_uart/uart0/tx_count16[2]~FF .SR_POLARITY = 1'b0;
    defparam \per_uart/uart0/tx_count16[2]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/tx_count16[2]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/tx_count16[2]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/tx_count16[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/tx_count16[3]~FF  (.D(\per_uart/uart0/n419 ), .CE(ceg_net203), 
           .CLK(\clk~O ), .SR(resetn), .Q(\per_uart/uart0/tx_count16[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(157)
    defparam \per_uart/uart0/tx_count16[3]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/tx_count16[3]~FF .CE_POLARITY = 1'b0;
    defparam \per_uart/uart0/tx_count16[3]~FF .SR_POLARITY = 1'b0;
    defparam \per_uart/uart0/tx_count16[3]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/tx_count16[3]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/tx_count16[3]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/tx_count16[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/txd_reg[1]~FF  (.D(\per_uart/uart0/n437 ), .CE(ceg_net159), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/uart0/txd_reg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(157)
    defparam \per_uart/uart0/txd_reg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/txd_reg[1]~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/uart0/txd_reg[1]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/uart0/txd_reg[1]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/txd_reg[1]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/txd_reg[1]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/txd_reg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/txd_reg[2]~FF  (.D(\per_uart/uart0/n436 ), .CE(ceg_net159), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/uart0/txd_reg[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(157)
    defparam \per_uart/uart0/txd_reg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/txd_reg[2]~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/uart0/txd_reg[2]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/uart0/txd_reg[2]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/txd_reg[2]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/txd_reg[2]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/txd_reg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/txd_reg[3]~FF  (.D(\per_uart/uart0/n435 ), .CE(ceg_net159), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/uart0/txd_reg[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(157)
    defparam \per_uart/uart0/txd_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/txd_reg[3]~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/uart0/txd_reg[3]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/uart0/txd_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/txd_reg[3]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/txd_reg[3]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/txd_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/txd_reg[4]~FF  (.D(\per_uart/uart0/n434 ), .CE(ceg_net159), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/uart0/txd_reg[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(157)
    defparam \per_uart/uart0/txd_reg[4]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/txd_reg[4]~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/uart0/txd_reg[4]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/uart0/txd_reg[4]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/txd_reg[4]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/txd_reg[4]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/txd_reg[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/txd_reg[5]~FF  (.D(\per_uart/uart0/n433 ), .CE(ceg_net159), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/uart0/txd_reg[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(157)
    defparam \per_uart/uart0/txd_reg[5]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/txd_reg[5]~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/uart0/txd_reg[5]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/uart0/txd_reg[5]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/txd_reg[5]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/txd_reg[5]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/txd_reg[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/txd_reg[6]~FF  (.D(\per_uart/uart0/n432 ), .CE(ceg_net159), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/uart0/txd_reg[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(157)
    defparam \per_uart/uart0/txd_reg[6]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/txd_reg[6]~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/uart0/txd_reg[6]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/uart0/txd_reg[6]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/txd_reg[6]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/txd_reg[6]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/txd_reg[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/txd_reg[7]~FF  (.D(\per_uart/uart0/n431 ), .CE(ceg_net159), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/uart0/txd_reg[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(157)
    defparam \per_uart/uart0/txd_reg[7]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/txd_reg[7]~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/uart0/txd_reg[7]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/uart0/txd_reg[7]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/txd_reg[7]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/txd_reg[7]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/txd_reg[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/tx_bitcount[1]~FF  (.D(\per_uart/uart0/n426 ), 
           .CE(ceg_net246), .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/uart0/tx_bitcount[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(157)
    defparam \per_uart/uart0/tx_bitcount[1]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/tx_bitcount[1]~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/uart0/tx_bitcount[1]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/uart0/tx_bitcount[1]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/tx_bitcount[1]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/tx_bitcount[1]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/tx_bitcount[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/tx_bitcount[2]~FF  (.D(\per_uart/uart0/n425 ), 
           .CE(ceg_net246), .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/uart0/tx_bitcount[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(157)
    defparam \per_uart/uart0/tx_bitcount[2]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/tx_bitcount[2]~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/uart0/tx_bitcount[2]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/uart0/tx_bitcount[2]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/tx_bitcount[2]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/tx_bitcount[2]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/tx_bitcount[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/tx_bitcount[3]~FF  (.D(\per_uart/uart0/n424 ), 
           .CE(ceg_net246), .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/uart0/tx_bitcount[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(157)
    defparam \per_uart/uart0/tx_bitcount[3]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/tx_bitcount[3]~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/uart0/tx_bitcount[3]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/uart0/tx_bitcount[3]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/tx_bitcount[3]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/tx_bitcount[3]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/tx_bitcount[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/enable16_counter[1]~FF  (.D(\per_uart/uart0/n732 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\per_uart/uart0/n552 ), .Q(\per_uart/uart0/enable16_counter[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(44)
    defparam \per_uart/uart0/enable16_counter[1]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/enable16_counter[1]~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/uart0/enable16_counter[1]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/uart0/enable16_counter[1]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/enable16_counter[1]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/enable16_counter[1]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/enable16_counter[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/enable16_counter[2]~FF  (.D(\per_uart/uart0/n737 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\per_uart/uart0/n552 ), .Q(\per_uart/uart0/enable16_counter[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(44)
    defparam \per_uart/uart0/enable16_counter[2]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/enable16_counter[2]~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/uart0/enable16_counter[2]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/uart0/enable16_counter[2]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/enable16_counter[2]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/enable16_counter[2]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/enable16_counter[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/enable16_counter[3]~FF  (.D(\per_uart/uart0/n742 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\per_uart/uart0/n552 ), .Q(\per_uart/uart0/enable16_counter[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(44)
    defparam \per_uart/uart0/enable16_counter[3]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/enable16_counter[3]~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/uart0/enable16_counter[3]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/uart0/enable16_counter[3]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/enable16_counter[3]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/enable16_counter[3]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/uart0/enable16_counter[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/uart0/enable16_counter[4]~FF  (.D(\per_uart/uart0/n747 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\per_uart/uart0/n552 ), .Q(\per_uart/uart0/enable16_counter[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/uart.v(44)
    defparam \per_uart/uart0/enable16_counter[4]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/uart0/enable16_counter[4]~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/uart0/enable16_counter[4]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/uart0/enable16_counter[4]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/uart0/enable16_counter[4]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/uart0/enable16_counter[4]~FF .SR_VALUE = 1'b1;
    defparam \per_uart/uart0/enable16_counter[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/d_in_uart[1]~FF  (.D(\mem_wdata[1] ), .CE(\per_uart/n15 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/d_in_uart[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/perip_uart.v(42)
    defparam \per_uart/d_in_uart[1]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/d_in_uart[1]~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/d_in_uart[1]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/d_in_uart[1]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/d_in_uart[1]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/d_in_uart[1]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/d_in_uart[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/d_in_uart[2]~FF  (.D(\mem_wdata[2] ), .CE(\per_uart/n15 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/d_in_uart[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/perip_uart.v(42)
    defparam \per_uart/d_in_uart[2]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/d_in_uart[2]~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/d_in_uart[2]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/d_in_uart[2]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/d_in_uart[2]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/d_in_uart[2]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/d_in_uart[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/d_in_uart[3]~FF  (.D(\mem_wdata[3] ), .CE(\per_uart/n15 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/d_in_uart[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/perip_uart.v(42)
    defparam \per_uart/d_in_uart[3]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/d_in_uart[3]~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/d_in_uart[3]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/d_in_uart[3]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/d_in_uart[3]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/d_in_uart[3]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/d_in_uart[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/d_in_uart[4]~FF  (.D(\mem_wdata[4] ), .CE(\per_uart/n15 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/d_in_uart[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/perip_uart.v(42)
    defparam \per_uart/d_in_uart[4]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/d_in_uart[4]~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/d_in_uart[4]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/d_in_uart[4]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/d_in_uart[4]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/d_in_uart[4]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/d_in_uart[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/d_in_uart[5]~FF  (.D(\mem_wdata[5] ), .CE(\per_uart/n15 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/d_in_uart[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/perip_uart.v(42)
    defparam \per_uart/d_in_uart[5]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/d_in_uart[5]~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/d_in_uart[5]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/d_in_uart[5]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/d_in_uart[5]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/d_in_uart[5]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/d_in_uart[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/d_in_uart[6]~FF  (.D(\mem_wdata[6] ), .CE(\per_uart/n15 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/d_in_uart[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/perip_uart.v(42)
    defparam \per_uart/d_in_uart[6]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/d_in_uart[6]~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/d_in_uart[6]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/d_in_uart[6]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/d_in_uart[6]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/d_in_uart[6]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/d_in_uart[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \per_uart/d_in_uart[7]~FF  (.D(\mem_wdata[7] ), .CE(\per_uart/n15 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\per_uart/d_in_uart[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/uart/perip_uart.v(42)
    defparam \per_uart/d_in_uart[7]~FF .CLK_POLARITY = 1'b1;
    defparam \per_uart/d_in_uart[7]~FF .CE_POLARITY = 1'b1;
    defparam \per_uart/d_in_uart[7]~FF .SR_POLARITY = 1'b1;
    defparam \per_uart/d_in_uart[7]~FF .D_POLARITY = 1'b1;
    defparam \per_uart/d_in_uart[7]~FF .SR_SYNC = 1'b1;
    defparam \per_uart/d_in_uart[7]~FF .SR_VALUE = 1'b0;
    defparam \per_uart/d_in_uart[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/A[0]~FF  (.D(\mem_wdata[0] ), .CE(\mult1/n402 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult1/A[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(53)
    defparam \mult1/A[0]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/A[0]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/A[0]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/A[0]~FF .D_POLARITY = 1'b1;
    defparam \mult1/A[0]~FF .SR_SYNC = 1'b1;
    defparam \mult1/A[0]~FF .SR_VALUE = 1'b0;
    defparam \mult1/A[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/B[0]~FF  (.D(\mem_wdata[0] ), .CE(\mult1/n403 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult1/B[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(53)
    defparam \mult1/B[0]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/B[0]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/B[0]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/B[0]~FF .D_POLARITY = 1'b1;
    defparam \mult1/B[0]~FF .SR_SYNC = 1'b1;
    defparam \mult1/B[0]~FF .SR_VALUE = 1'b0;
    defparam \mult1/B[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult_dout[0]~FF  (.D(\mult1/n201 ), .CE(\mult1/n165 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult_dout[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(65)
    defparam \mult_dout[0]~FF .CLK_POLARITY = 1'b1;
    defparam \mult_dout[0]~FF .CE_POLARITY = 1'b1;
    defparam \mult_dout[0]~FF .SR_POLARITY = 1'b0;
    defparam \mult_dout[0]~FF .D_POLARITY = 1'b1;
    defparam \mult_dout[0]~FF .SR_SYNC = 1'b1;
    defparam \mult_dout[0]~FF .SR_VALUE = 1'b0;
    defparam \mult_dout[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/init~FF  (.D(\mem_wdata[0] ), .CE(\mult1/n404 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult1/init )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(53)
    defparam \mult1/init~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/init~FF .CE_POLARITY = 1'b1;
    defparam \mult1/init~FF .SR_POLARITY = 1'b0;
    defparam \mult1/init~FF .D_POLARITY = 1'b1;
    defparam \mult1/init~FF .SR_SYNC = 1'b1;
    defparam \mult1/init~FF .SR_VALUE = 1'b0;
    defparam \mult1/init~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/A[1]~FF  (.D(\mem_wdata[1] ), .CE(\mult1/n402 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult1/A[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(53)
    defparam \mult1/A[1]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/A[1]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/A[1]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/A[1]~FF .D_POLARITY = 1'b1;
    defparam \mult1/A[1]~FF .SR_SYNC = 1'b1;
    defparam \mult1/A[1]~FF .SR_VALUE = 1'b0;
    defparam \mult1/A[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/A[2]~FF  (.D(\mem_wdata[2] ), .CE(\mult1/n402 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult1/A[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(53)
    defparam \mult1/A[2]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/A[2]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/A[2]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/A[2]~FF .D_POLARITY = 1'b1;
    defparam \mult1/A[2]~FF .SR_SYNC = 1'b1;
    defparam \mult1/A[2]~FF .SR_VALUE = 1'b0;
    defparam \mult1/A[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/A[3]~FF  (.D(\mem_wdata[3] ), .CE(\mult1/n402 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult1/A[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(53)
    defparam \mult1/A[3]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/A[3]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/A[3]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/A[3]~FF .D_POLARITY = 1'b1;
    defparam \mult1/A[3]~FF .SR_SYNC = 1'b1;
    defparam \mult1/A[3]~FF .SR_VALUE = 1'b0;
    defparam \mult1/A[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/A[4]~FF  (.D(\mem_wdata[4] ), .CE(\mult1/n402 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult1/A[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(53)
    defparam \mult1/A[4]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/A[4]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/A[4]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/A[4]~FF .D_POLARITY = 1'b1;
    defparam \mult1/A[4]~FF .SR_SYNC = 1'b1;
    defparam \mult1/A[4]~FF .SR_VALUE = 1'b0;
    defparam \mult1/A[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/A[5]~FF  (.D(\mem_wdata[5] ), .CE(\mult1/n402 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult1/A[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(53)
    defparam \mult1/A[5]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/A[5]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/A[5]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/A[5]~FF .D_POLARITY = 1'b1;
    defparam \mult1/A[5]~FF .SR_SYNC = 1'b1;
    defparam \mult1/A[5]~FF .SR_VALUE = 1'b0;
    defparam \mult1/A[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/A[6]~FF  (.D(\mem_wdata[6] ), .CE(\mult1/n402 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult1/A[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(53)
    defparam \mult1/A[6]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/A[6]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/A[6]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/A[6]~FF .D_POLARITY = 1'b1;
    defparam \mult1/A[6]~FF .SR_SYNC = 1'b1;
    defparam \mult1/A[6]~FF .SR_VALUE = 1'b0;
    defparam \mult1/A[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/A[7]~FF  (.D(\mem_wdata[7] ), .CE(\mult1/n402 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult1/A[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(53)
    defparam \mult1/A[7]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/A[7]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/A[7]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/A[7]~FF .D_POLARITY = 1'b1;
    defparam \mult1/A[7]~FF .SR_SYNC = 1'b1;
    defparam \mult1/A[7]~FF .SR_VALUE = 1'b0;
    defparam \mult1/A[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/A[8]~FF  (.D(\mem_wdata[8] ), .CE(\mult1/n402 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult1/A[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(53)
    defparam \mult1/A[8]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/A[8]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/A[8]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/A[8]~FF .D_POLARITY = 1'b1;
    defparam \mult1/A[8]~FF .SR_SYNC = 1'b1;
    defparam \mult1/A[8]~FF .SR_VALUE = 1'b0;
    defparam \mult1/A[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/A[9]~FF  (.D(\mem_wdata[9] ), .CE(\mult1/n402 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult1/A[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(53)
    defparam \mult1/A[9]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/A[9]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/A[9]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/A[9]~FF .D_POLARITY = 1'b1;
    defparam \mult1/A[9]~FF .SR_SYNC = 1'b1;
    defparam \mult1/A[9]~FF .SR_VALUE = 1'b0;
    defparam \mult1/A[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/A[10]~FF  (.D(\mem_wdata[10] ), .CE(\mult1/n402 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult1/A[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(53)
    defparam \mult1/A[10]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/A[10]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/A[10]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/A[10]~FF .D_POLARITY = 1'b1;
    defparam \mult1/A[10]~FF .SR_SYNC = 1'b1;
    defparam \mult1/A[10]~FF .SR_VALUE = 1'b0;
    defparam \mult1/A[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/A[11]~FF  (.D(\mem_wdata[11] ), .CE(\mult1/n402 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult1/A[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(53)
    defparam \mult1/A[11]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/A[11]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/A[11]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/A[11]~FF .D_POLARITY = 1'b1;
    defparam \mult1/A[11]~FF .SR_SYNC = 1'b1;
    defparam \mult1/A[11]~FF .SR_VALUE = 1'b0;
    defparam \mult1/A[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/A[12]~FF  (.D(\mem_wdata[12] ), .CE(\mult1/n402 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult1/A[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(53)
    defparam \mult1/A[12]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/A[12]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/A[12]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/A[12]~FF .D_POLARITY = 1'b1;
    defparam \mult1/A[12]~FF .SR_SYNC = 1'b1;
    defparam \mult1/A[12]~FF .SR_VALUE = 1'b0;
    defparam \mult1/A[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/A[13]~FF  (.D(\mem_wdata[13] ), .CE(\mult1/n402 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult1/A[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(53)
    defparam \mult1/A[13]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/A[13]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/A[13]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/A[13]~FF .D_POLARITY = 1'b1;
    defparam \mult1/A[13]~FF .SR_SYNC = 1'b1;
    defparam \mult1/A[13]~FF .SR_VALUE = 1'b0;
    defparam \mult1/A[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/A[14]~FF  (.D(\mem_wdata[14] ), .CE(\mult1/n402 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult1/A[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(53)
    defparam \mult1/A[14]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/A[14]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/A[14]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/A[14]~FF .D_POLARITY = 1'b1;
    defparam \mult1/A[14]~FF .SR_SYNC = 1'b1;
    defparam \mult1/A[14]~FF .SR_VALUE = 1'b0;
    defparam \mult1/A[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/A[15]~FF  (.D(\mem_wdata[15] ), .CE(\mult1/n402 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult1/A[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(53)
    defparam \mult1/A[15]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/A[15]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/A[15]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/A[15]~FF .D_POLARITY = 1'b1;
    defparam \mult1/A[15]~FF .SR_SYNC = 1'b1;
    defparam \mult1/A[15]~FF .SR_VALUE = 1'b0;
    defparam \mult1/A[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/B[1]~FF  (.D(\mem_wdata[1] ), .CE(\mult1/n403 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult1/B[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(53)
    defparam \mult1/B[1]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/B[1]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/B[1]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/B[1]~FF .D_POLARITY = 1'b1;
    defparam \mult1/B[1]~FF .SR_SYNC = 1'b1;
    defparam \mult1/B[1]~FF .SR_VALUE = 1'b0;
    defparam \mult1/B[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/B[2]~FF  (.D(\mem_wdata[2] ), .CE(\mult1/n403 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult1/B[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(53)
    defparam \mult1/B[2]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/B[2]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/B[2]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/B[2]~FF .D_POLARITY = 1'b1;
    defparam \mult1/B[2]~FF .SR_SYNC = 1'b1;
    defparam \mult1/B[2]~FF .SR_VALUE = 1'b0;
    defparam \mult1/B[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/B[3]~FF  (.D(\mem_wdata[3] ), .CE(\mult1/n403 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult1/B[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(53)
    defparam \mult1/B[3]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/B[3]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/B[3]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/B[3]~FF .D_POLARITY = 1'b1;
    defparam \mult1/B[3]~FF .SR_SYNC = 1'b1;
    defparam \mult1/B[3]~FF .SR_VALUE = 1'b0;
    defparam \mult1/B[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/B[4]~FF  (.D(\mem_wdata[4] ), .CE(\mult1/n403 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult1/B[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(53)
    defparam \mult1/B[4]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/B[4]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/B[4]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/B[4]~FF .D_POLARITY = 1'b1;
    defparam \mult1/B[4]~FF .SR_SYNC = 1'b1;
    defparam \mult1/B[4]~FF .SR_VALUE = 1'b0;
    defparam \mult1/B[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/B[5]~FF  (.D(\mem_wdata[5] ), .CE(\mult1/n403 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult1/B[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(53)
    defparam \mult1/B[5]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/B[5]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/B[5]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/B[5]~FF .D_POLARITY = 1'b1;
    defparam \mult1/B[5]~FF .SR_SYNC = 1'b1;
    defparam \mult1/B[5]~FF .SR_VALUE = 1'b0;
    defparam \mult1/B[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/B[6]~FF  (.D(\mem_wdata[6] ), .CE(\mult1/n403 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult1/B[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(53)
    defparam \mult1/B[6]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/B[6]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/B[6]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/B[6]~FF .D_POLARITY = 1'b1;
    defparam \mult1/B[6]~FF .SR_SYNC = 1'b1;
    defparam \mult1/B[6]~FF .SR_VALUE = 1'b0;
    defparam \mult1/B[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/B[7]~FF  (.D(\mem_wdata[7] ), .CE(\mult1/n403 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult1/B[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(53)
    defparam \mult1/B[7]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/B[7]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/B[7]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/B[7]~FF .D_POLARITY = 1'b1;
    defparam \mult1/B[7]~FF .SR_SYNC = 1'b1;
    defparam \mult1/B[7]~FF .SR_VALUE = 1'b0;
    defparam \mult1/B[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/B[8]~FF  (.D(\mem_wdata[8] ), .CE(\mult1/n403 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult1/B[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(53)
    defparam \mult1/B[8]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/B[8]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/B[8]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/B[8]~FF .D_POLARITY = 1'b1;
    defparam \mult1/B[8]~FF .SR_SYNC = 1'b1;
    defparam \mult1/B[8]~FF .SR_VALUE = 1'b0;
    defparam \mult1/B[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/B[9]~FF  (.D(\mem_wdata[9] ), .CE(\mult1/n403 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult1/B[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(53)
    defparam \mult1/B[9]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/B[9]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/B[9]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/B[9]~FF .D_POLARITY = 1'b1;
    defparam \mult1/B[9]~FF .SR_SYNC = 1'b1;
    defparam \mult1/B[9]~FF .SR_VALUE = 1'b0;
    defparam \mult1/B[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/B[10]~FF  (.D(\mem_wdata[10] ), .CE(\mult1/n403 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult1/B[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(53)
    defparam \mult1/B[10]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/B[10]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/B[10]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/B[10]~FF .D_POLARITY = 1'b1;
    defparam \mult1/B[10]~FF .SR_SYNC = 1'b1;
    defparam \mult1/B[10]~FF .SR_VALUE = 1'b0;
    defparam \mult1/B[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/B[11]~FF  (.D(\mem_wdata[11] ), .CE(\mult1/n403 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult1/B[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(53)
    defparam \mult1/B[11]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/B[11]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/B[11]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/B[11]~FF .D_POLARITY = 1'b1;
    defparam \mult1/B[11]~FF .SR_SYNC = 1'b1;
    defparam \mult1/B[11]~FF .SR_VALUE = 1'b0;
    defparam \mult1/B[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/B[12]~FF  (.D(\mem_wdata[12] ), .CE(\mult1/n403 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult1/B[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(53)
    defparam \mult1/B[12]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/B[12]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/B[12]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/B[12]~FF .D_POLARITY = 1'b1;
    defparam \mult1/B[12]~FF .SR_SYNC = 1'b1;
    defparam \mult1/B[12]~FF .SR_VALUE = 1'b0;
    defparam \mult1/B[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/B[13]~FF  (.D(\mem_wdata[13] ), .CE(\mult1/n403 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult1/B[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(53)
    defparam \mult1/B[13]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/B[13]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/B[13]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/B[13]~FF .D_POLARITY = 1'b1;
    defparam \mult1/B[13]~FF .SR_SYNC = 1'b1;
    defparam \mult1/B[13]~FF .SR_VALUE = 1'b0;
    defparam \mult1/B[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/B[14]~FF  (.D(\mem_wdata[14] ), .CE(\mult1/n403 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult1/B[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(53)
    defparam \mult1/B[14]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/B[14]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/B[14]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/B[14]~FF .D_POLARITY = 1'b1;
    defparam \mult1/B[14]~FF .SR_SYNC = 1'b1;
    defparam \mult1/B[14]~FF .SR_VALUE = 1'b0;
    defparam \mult1/B[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/B[15]~FF  (.D(\mem_wdata[15] ), .CE(\mult1/n403 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult1/B[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(53)
    defparam \mult1/B[15]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/B[15]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/B[15]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/B[15]~FF .D_POLARITY = 1'b1;
    defparam \mult1/B[15]~FF .SR_SYNC = 1'b1;
    defparam \mult1/B[15]~FF .SR_VALUE = 1'b0;
    defparam \mult1/B[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult_dout[1]~FF  (.D(\mult1/n200 ), .CE(\mult1/n165 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult_dout[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(65)
    defparam \mult_dout[1]~FF .CLK_POLARITY = 1'b1;
    defparam \mult_dout[1]~FF .CE_POLARITY = 1'b1;
    defparam \mult_dout[1]~FF .SR_POLARITY = 1'b0;
    defparam \mult_dout[1]~FF .D_POLARITY = 1'b1;
    defparam \mult_dout[1]~FF .SR_SYNC = 1'b1;
    defparam \mult_dout[1]~FF .SR_VALUE = 1'b0;
    defparam \mult_dout[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult_dout[2]~FF  (.D(\mult1/n199 ), .CE(\mult1/n165 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult_dout[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(65)
    defparam \mult_dout[2]~FF .CLK_POLARITY = 1'b1;
    defparam \mult_dout[2]~FF .CE_POLARITY = 1'b1;
    defparam \mult_dout[2]~FF .SR_POLARITY = 1'b0;
    defparam \mult_dout[2]~FF .D_POLARITY = 1'b1;
    defparam \mult_dout[2]~FF .SR_SYNC = 1'b1;
    defparam \mult_dout[2]~FF .SR_VALUE = 1'b0;
    defparam \mult_dout[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult_dout[3]~FF  (.D(\mult1/n198 ), .CE(\mult1/n165 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult_dout[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(65)
    defparam \mult_dout[3]~FF .CLK_POLARITY = 1'b1;
    defparam \mult_dout[3]~FF .CE_POLARITY = 1'b1;
    defparam \mult_dout[3]~FF .SR_POLARITY = 1'b0;
    defparam \mult_dout[3]~FF .D_POLARITY = 1'b1;
    defparam \mult_dout[3]~FF .SR_SYNC = 1'b1;
    defparam \mult_dout[3]~FF .SR_VALUE = 1'b0;
    defparam \mult_dout[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult_dout[4]~FF  (.D(\mult1/n197 ), .CE(\mult1/n165 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult_dout[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(65)
    defparam \mult_dout[4]~FF .CLK_POLARITY = 1'b1;
    defparam \mult_dout[4]~FF .CE_POLARITY = 1'b1;
    defparam \mult_dout[4]~FF .SR_POLARITY = 1'b0;
    defparam \mult_dout[4]~FF .D_POLARITY = 1'b1;
    defparam \mult_dout[4]~FF .SR_SYNC = 1'b1;
    defparam \mult_dout[4]~FF .SR_VALUE = 1'b0;
    defparam \mult_dout[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult_dout[5]~FF  (.D(\mult1/n196 ), .CE(\mult1/n165 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult_dout[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(65)
    defparam \mult_dout[5]~FF .CLK_POLARITY = 1'b1;
    defparam \mult_dout[5]~FF .CE_POLARITY = 1'b1;
    defparam \mult_dout[5]~FF .SR_POLARITY = 1'b0;
    defparam \mult_dout[5]~FF .D_POLARITY = 1'b1;
    defparam \mult_dout[5]~FF .SR_SYNC = 1'b1;
    defparam \mult_dout[5]~FF .SR_VALUE = 1'b0;
    defparam \mult_dout[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult_dout[6]~FF  (.D(\mult1/n195 ), .CE(\mult1/n165 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult_dout[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(65)
    defparam \mult_dout[6]~FF .CLK_POLARITY = 1'b1;
    defparam \mult_dout[6]~FF .CE_POLARITY = 1'b1;
    defparam \mult_dout[6]~FF .SR_POLARITY = 1'b0;
    defparam \mult_dout[6]~FF .D_POLARITY = 1'b1;
    defparam \mult_dout[6]~FF .SR_SYNC = 1'b1;
    defparam \mult_dout[6]~FF .SR_VALUE = 1'b0;
    defparam \mult_dout[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult_dout[7]~FF  (.D(\mult1/n194 ), .CE(\mult1/n165 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult_dout[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(65)
    defparam \mult_dout[7]~FF .CLK_POLARITY = 1'b1;
    defparam \mult_dout[7]~FF .CE_POLARITY = 1'b1;
    defparam \mult_dout[7]~FF .SR_POLARITY = 1'b0;
    defparam \mult_dout[7]~FF .D_POLARITY = 1'b1;
    defparam \mult_dout[7]~FF .SR_SYNC = 1'b1;
    defparam \mult_dout[7]~FF .SR_VALUE = 1'b0;
    defparam \mult_dout[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult_dout[8]~FF  (.D(\mult1/n193 ), .CE(\mult1/n165 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult_dout[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(65)
    defparam \mult_dout[8]~FF .CLK_POLARITY = 1'b1;
    defparam \mult_dout[8]~FF .CE_POLARITY = 1'b1;
    defparam \mult_dout[8]~FF .SR_POLARITY = 1'b0;
    defparam \mult_dout[8]~FF .D_POLARITY = 1'b1;
    defparam \mult_dout[8]~FF .SR_SYNC = 1'b1;
    defparam \mult_dout[8]~FF .SR_VALUE = 1'b0;
    defparam \mult_dout[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult_dout[9]~FF  (.D(\mult1/n192 ), .CE(\mult1/n165 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult_dout[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(65)
    defparam \mult_dout[9]~FF .CLK_POLARITY = 1'b1;
    defparam \mult_dout[9]~FF .CE_POLARITY = 1'b1;
    defparam \mult_dout[9]~FF .SR_POLARITY = 1'b0;
    defparam \mult_dout[9]~FF .D_POLARITY = 1'b1;
    defparam \mult_dout[9]~FF .SR_SYNC = 1'b1;
    defparam \mult_dout[9]~FF .SR_VALUE = 1'b0;
    defparam \mult_dout[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult_dout[10]~FF  (.D(\mult1/n191 ), .CE(\mult1/n165 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult_dout[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(65)
    defparam \mult_dout[10]~FF .CLK_POLARITY = 1'b1;
    defparam \mult_dout[10]~FF .CE_POLARITY = 1'b1;
    defparam \mult_dout[10]~FF .SR_POLARITY = 1'b0;
    defparam \mult_dout[10]~FF .D_POLARITY = 1'b1;
    defparam \mult_dout[10]~FF .SR_SYNC = 1'b1;
    defparam \mult_dout[10]~FF .SR_VALUE = 1'b0;
    defparam \mult_dout[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult_dout[11]~FF  (.D(\mult1/n190 ), .CE(\mult1/n165 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult_dout[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(65)
    defparam \mult_dout[11]~FF .CLK_POLARITY = 1'b1;
    defparam \mult_dout[11]~FF .CE_POLARITY = 1'b1;
    defparam \mult_dout[11]~FF .SR_POLARITY = 1'b0;
    defparam \mult_dout[11]~FF .D_POLARITY = 1'b1;
    defparam \mult_dout[11]~FF .SR_SYNC = 1'b1;
    defparam \mult_dout[11]~FF .SR_VALUE = 1'b0;
    defparam \mult_dout[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult_dout[12]~FF  (.D(\mult1/n189 ), .CE(\mult1/n165 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult_dout[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(65)
    defparam \mult_dout[12]~FF .CLK_POLARITY = 1'b1;
    defparam \mult_dout[12]~FF .CE_POLARITY = 1'b1;
    defparam \mult_dout[12]~FF .SR_POLARITY = 1'b0;
    defparam \mult_dout[12]~FF .D_POLARITY = 1'b1;
    defparam \mult_dout[12]~FF .SR_SYNC = 1'b1;
    defparam \mult_dout[12]~FF .SR_VALUE = 1'b0;
    defparam \mult_dout[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult_dout[13]~FF  (.D(\mult1/n188 ), .CE(\mult1/n165 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult_dout[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(65)
    defparam \mult_dout[13]~FF .CLK_POLARITY = 1'b1;
    defparam \mult_dout[13]~FF .CE_POLARITY = 1'b1;
    defparam \mult_dout[13]~FF .SR_POLARITY = 1'b0;
    defparam \mult_dout[13]~FF .D_POLARITY = 1'b1;
    defparam \mult_dout[13]~FF .SR_SYNC = 1'b1;
    defparam \mult_dout[13]~FF .SR_VALUE = 1'b0;
    defparam \mult_dout[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult_dout[14]~FF  (.D(\mult1/n187 ), .CE(\mult1/n165 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult_dout[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(65)
    defparam \mult_dout[14]~FF .CLK_POLARITY = 1'b1;
    defparam \mult_dout[14]~FF .CE_POLARITY = 1'b1;
    defparam \mult_dout[14]~FF .SR_POLARITY = 1'b0;
    defparam \mult_dout[14]~FF .D_POLARITY = 1'b1;
    defparam \mult_dout[14]~FF .SR_SYNC = 1'b1;
    defparam \mult_dout[14]~FF .SR_VALUE = 1'b0;
    defparam \mult_dout[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult_dout[15]~FF  (.D(\mult1/n186 ), .CE(\mult1/n165 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult_dout[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(65)
    defparam \mult_dout[15]~FF .CLK_POLARITY = 1'b1;
    defparam \mult_dout[15]~FF .CE_POLARITY = 1'b1;
    defparam \mult_dout[15]~FF .SR_POLARITY = 1'b0;
    defparam \mult_dout[15]~FF .D_POLARITY = 1'b1;
    defparam \mult_dout[15]~FF .SR_SYNC = 1'b1;
    defparam \mult_dout[15]~FF .SR_VALUE = 1'b0;
    defparam \mult_dout[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult_dout[16]~FF  (.D(\mult1/n185 ), .CE(\mult1/n165 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult_dout[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(65)
    defparam \mult_dout[16]~FF .CLK_POLARITY = 1'b1;
    defparam \mult_dout[16]~FF .CE_POLARITY = 1'b1;
    defparam \mult_dout[16]~FF .SR_POLARITY = 1'b0;
    defparam \mult_dout[16]~FF .D_POLARITY = 1'b1;
    defparam \mult_dout[16]~FF .SR_SYNC = 1'b1;
    defparam \mult_dout[16]~FF .SR_VALUE = 1'b0;
    defparam \mult_dout[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult_dout[17]~FF  (.D(\mult1/n184 ), .CE(\mult1/n165 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult_dout[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(65)
    defparam \mult_dout[17]~FF .CLK_POLARITY = 1'b1;
    defparam \mult_dout[17]~FF .CE_POLARITY = 1'b1;
    defparam \mult_dout[17]~FF .SR_POLARITY = 1'b0;
    defparam \mult_dout[17]~FF .D_POLARITY = 1'b1;
    defparam \mult_dout[17]~FF .SR_SYNC = 1'b1;
    defparam \mult_dout[17]~FF .SR_VALUE = 1'b0;
    defparam \mult_dout[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult_dout[18]~FF  (.D(\mult1/n183 ), .CE(\mult1/n165 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult_dout[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(65)
    defparam \mult_dout[18]~FF .CLK_POLARITY = 1'b1;
    defparam \mult_dout[18]~FF .CE_POLARITY = 1'b1;
    defparam \mult_dout[18]~FF .SR_POLARITY = 1'b0;
    defparam \mult_dout[18]~FF .D_POLARITY = 1'b1;
    defparam \mult_dout[18]~FF .SR_SYNC = 1'b1;
    defparam \mult_dout[18]~FF .SR_VALUE = 1'b0;
    defparam \mult_dout[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult_dout[19]~FF  (.D(\mult1/n182 ), .CE(\mult1/n165 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult_dout[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(65)
    defparam \mult_dout[19]~FF .CLK_POLARITY = 1'b1;
    defparam \mult_dout[19]~FF .CE_POLARITY = 1'b1;
    defparam \mult_dout[19]~FF .SR_POLARITY = 1'b0;
    defparam \mult_dout[19]~FF .D_POLARITY = 1'b1;
    defparam \mult_dout[19]~FF .SR_SYNC = 1'b1;
    defparam \mult_dout[19]~FF .SR_VALUE = 1'b0;
    defparam \mult_dout[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult_dout[20]~FF  (.D(\mult1/n181 ), .CE(\mult1/n165 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult_dout[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(65)
    defparam \mult_dout[20]~FF .CLK_POLARITY = 1'b1;
    defparam \mult_dout[20]~FF .CE_POLARITY = 1'b1;
    defparam \mult_dout[20]~FF .SR_POLARITY = 1'b0;
    defparam \mult_dout[20]~FF .D_POLARITY = 1'b1;
    defparam \mult_dout[20]~FF .SR_SYNC = 1'b1;
    defparam \mult_dout[20]~FF .SR_VALUE = 1'b0;
    defparam \mult_dout[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult_dout[21]~FF  (.D(\mult1/n180 ), .CE(\mult1/n165 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult_dout[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(65)
    defparam \mult_dout[21]~FF .CLK_POLARITY = 1'b1;
    defparam \mult_dout[21]~FF .CE_POLARITY = 1'b1;
    defparam \mult_dout[21]~FF .SR_POLARITY = 1'b0;
    defparam \mult_dout[21]~FF .D_POLARITY = 1'b1;
    defparam \mult_dout[21]~FF .SR_SYNC = 1'b1;
    defparam \mult_dout[21]~FF .SR_VALUE = 1'b0;
    defparam \mult_dout[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult_dout[22]~FF  (.D(\mult1/n179 ), .CE(\mult1/n165 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult_dout[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(65)
    defparam \mult_dout[22]~FF .CLK_POLARITY = 1'b1;
    defparam \mult_dout[22]~FF .CE_POLARITY = 1'b1;
    defparam \mult_dout[22]~FF .SR_POLARITY = 1'b0;
    defparam \mult_dout[22]~FF .D_POLARITY = 1'b1;
    defparam \mult_dout[22]~FF .SR_SYNC = 1'b1;
    defparam \mult_dout[22]~FF .SR_VALUE = 1'b0;
    defparam \mult_dout[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult_dout[23]~FF  (.D(\mult1/n178 ), .CE(\mult1/n165 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult_dout[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(65)
    defparam \mult_dout[23]~FF .CLK_POLARITY = 1'b1;
    defparam \mult_dout[23]~FF .CE_POLARITY = 1'b1;
    defparam \mult_dout[23]~FF .SR_POLARITY = 1'b0;
    defparam \mult_dout[23]~FF .D_POLARITY = 1'b1;
    defparam \mult_dout[23]~FF .SR_SYNC = 1'b1;
    defparam \mult_dout[23]~FF .SR_VALUE = 1'b0;
    defparam \mult_dout[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult_dout[24]~FF  (.D(\mult1/n177 ), .CE(\mult1/n165 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult_dout[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(65)
    defparam \mult_dout[24]~FF .CLK_POLARITY = 1'b1;
    defparam \mult_dout[24]~FF .CE_POLARITY = 1'b1;
    defparam \mult_dout[24]~FF .SR_POLARITY = 1'b0;
    defparam \mult_dout[24]~FF .D_POLARITY = 1'b1;
    defparam \mult_dout[24]~FF .SR_SYNC = 1'b1;
    defparam \mult_dout[24]~FF .SR_VALUE = 1'b0;
    defparam \mult_dout[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult_dout[25]~FF  (.D(\mult1/n176 ), .CE(\mult1/n165 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult_dout[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(65)
    defparam \mult_dout[25]~FF .CLK_POLARITY = 1'b1;
    defparam \mult_dout[25]~FF .CE_POLARITY = 1'b1;
    defparam \mult_dout[25]~FF .SR_POLARITY = 1'b0;
    defparam \mult_dout[25]~FF .D_POLARITY = 1'b1;
    defparam \mult_dout[25]~FF .SR_SYNC = 1'b1;
    defparam \mult_dout[25]~FF .SR_VALUE = 1'b0;
    defparam \mult_dout[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult_dout[26]~FF  (.D(\mult1/n175 ), .CE(\mult1/n165 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult_dout[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(65)
    defparam \mult_dout[26]~FF .CLK_POLARITY = 1'b1;
    defparam \mult_dout[26]~FF .CE_POLARITY = 1'b1;
    defparam \mult_dout[26]~FF .SR_POLARITY = 1'b0;
    defparam \mult_dout[26]~FF .D_POLARITY = 1'b1;
    defparam \mult_dout[26]~FF .SR_SYNC = 1'b1;
    defparam \mult_dout[26]~FF .SR_VALUE = 1'b0;
    defparam \mult_dout[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult_dout[27]~FF  (.D(\mult1/n174 ), .CE(\mult1/n165 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult_dout[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(65)
    defparam \mult_dout[27]~FF .CLK_POLARITY = 1'b1;
    defparam \mult_dout[27]~FF .CE_POLARITY = 1'b1;
    defparam \mult_dout[27]~FF .SR_POLARITY = 1'b0;
    defparam \mult_dout[27]~FF .D_POLARITY = 1'b1;
    defparam \mult_dout[27]~FF .SR_SYNC = 1'b1;
    defparam \mult_dout[27]~FF .SR_VALUE = 1'b0;
    defparam \mult_dout[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult_dout[28]~FF  (.D(\mult1/n173 ), .CE(\mult1/n165 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult_dout[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(65)
    defparam \mult_dout[28]~FF .CLK_POLARITY = 1'b1;
    defparam \mult_dout[28]~FF .CE_POLARITY = 1'b1;
    defparam \mult_dout[28]~FF .SR_POLARITY = 1'b0;
    defparam \mult_dout[28]~FF .D_POLARITY = 1'b1;
    defparam \mult_dout[28]~FF .SR_SYNC = 1'b1;
    defparam \mult_dout[28]~FF .SR_VALUE = 1'b0;
    defparam \mult_dout[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult_dout[29]~FF  (.D(\mult1/n172 ), .CE(\mult1/n165 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult_dout[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(65)
    defparam \mult_dout[29]~FF .CLK_POLARITY = 1'b1;
    defparam \mult_dout[29]~FF .CE_POLARITY = 1'b1;
    defparam \mult_dout[29]~FF .SR_POLARITY = 1'b0;
    defparam \mult_dout[29]~FF .D_POLARITY = 1'b1;
    defparam \mult_dout[29]~FF .SR_SYNC = 1'b1;
    defparam \mult_dout[29]~FF .SR_VALUE = 1'b0;
    defparam \mult_dout[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult_dout[30]~FF  (.D(\mult1/n171 ), .CE(\mult1/n165 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult_dout[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(65)
    defparam \mult_dout[30]~FF .CLK_POLARITY = 1'b1;
    defparam \mult_dout[30]~FF .CE_POLARITY = 1'b1;
    defparam \mult_dout[30]~FF .SR_POLARITY = 1'b0;
    defparam \mult_dout[30]~FF .D_POLARITY = 1'b1;
    defparam \mult_dout[30]~FF .SR_SYNC = 1'b1;
    defparam \mult_dout[30]~FF .SR_VALUE = 1'b0;
    defparam \mult_dout[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult_dout[31]~FF  (.D(\mult1/n170 ), .CE(\mult1/n165 ), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult_dout[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/perip_mult.v(65)
    defparam \mult_dout[31]~FF .CLK_POLARITY = 1'b1;
    defparam \mult_dout[31]~FF .CE_POLARITY = 1'b1;
    defparam \mult_dout[31]~FF .SR_POLARITY = 1'b0;
    defparam \mult_dout[31]~FF .D_POLARITY = 1'b1;
    defparam \mult_dout[31]~FF .SR_SYNC = 1'b1;
    defparam \mult_dout[31]~FF .SR_VALUE = 1'b0;
    defparam \mult_dout[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/result[0]~FF  (.D(\mult1/mult1/n132 ), .CE(ceg_net913), 
           .CLK(\clk~O ), .SR(resetn), .Q(\mult1/result[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/result[0]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/result[0]~FF .CE_POLARITY = 1'b0;
    defparam \mult1/result[0]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/result[0]~FF .D_POLARITY = 1'b1;
    defparam \mult1/result[0]~FF .SR_SYNC = 1'b0;
    defparam \mult1/result[0]~FF .SR_VALUE = 1'b0;
    defparam \mult1/result[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/state[0]~FF  (.D(\mult1/mult1/n64 ), .CE(ceg_net252), 
           .CLK(\clk~O ), .SR(resetn), .Q(\mult1/mult1/state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/state[0]~FF .CE_POLARITY = 1'b0;
    defparam \mult1/mult1/state[0]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/mult1/state[0]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/state[0]~FF .SR_SYNC = 1'b0;
    defparam \mult1/mult1/state[0]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/A[0]~FF  (.D(\mult1/mult1/n81 ), .CE(ceg_net839), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/A[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/A[0]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/A[0]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/A[0]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/A[0]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/A[0]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/A[0]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/A[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/B[0]~FF  (.D(\mult1/mult1/n98 ), .CE(ceg_net839), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/B[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/B[0]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/B[0]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/B[0]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/B[0]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/B[0]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/B[0]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/B[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/count[0]~FF  (.D(\mult1/mult1/n138 ), .CE(ceg_net847), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/count[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/count[0]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/count[0]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/count[0]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/count[0]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/count[0]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/count[0]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/count[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/done~FF  (.D(\mult1/mult1/n99 ), .CE(ceg_net564), .CLK(\clk~O ), 
           .SR(resetn), .Q(\mult1/done )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/done~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/done~FF .CE_POLARITY = 1'b0;
    defparam \mult1/done~FF .SR_POLARITY = 1'b0;
    defparam \mult1/done~FF .D_POLARITY = 1'b1;
    defparam \mult1/done~FF .SR_SYNC = 1'b0;
    defparam \mult1/done~FF .SR_VALUE = 1'b0;
    defparam \mult1/done~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/result[1]~FF  (.D(\mult1/mult1/n131 ), .CE(ceg_net913), 
           .CLK(\clk~O ), .SR(resetn), .Q(\mult1/result[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/result[1]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/result[1]~FF .CE_POLARITY = 1'b0;
    defparam \mult1/result[1]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/result[1]~FF .D_POLARITY = 1'b1;
    defparam \mult1/result[1]~FF .SR_SYNC = 1'b0;
    defparam \mult1/result[1]~FF .SR_VALUE = 1'b0;
    defparam \mult1/result[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/result[2]~FF  (.D(\mult1/mult1/n130 ), .CE(ceg_net913), 
           .CLK(\clk~O ), .SR(resetn), .Q(\mult1/result[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/result[2]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/result[2]~FF .CE_POLARITY = 1'b0;
    defparam \mult1/result[2]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/result[2]~FF .D_POLARITY = 1'b1;
    defparam \mult1/result[2]~FF .SR_SYNC = 1'b0;
    defparam \mult1/result[2]~FF .SR_VALUE = 1'b0;
    defparam \mult1/result[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/result[3]~FF  (.D(\mult1/mult1/n129 ), .CE(ceg_net913), 
           .CLK(\clk~O ), .SR(resetn), .Q(\mult1/result[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/result[3]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/result[3]~FF .CE_POLARITY = 1'b0;
    defparam \mult1/result[3]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/result[3]~FF .D_POLARITY = 1'b1;
    defparam \mult1/result[3]~FF .SR_SYNC = 1'b0;
    defparam \mult1/result[3]~FF .SR_VALUE = 1'b0;
    defparam \mult1/result[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/result[4]~FF  (.D(\mult1/mult1/n128 ), .CE(ceg_net913), 
           .CLK(\clk~O ), .SR(resetn), .Q(\mult1/result[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/result[4]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/result[4]~FF .CE_POLARITY = 1'b0;
    defparam \mult1/result[4]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/result[4]~FF .D_POLARITY = 1'b1;
    defparam \mult1/result[4]~FF .SR_SYNC = 1'b0;
    defparam \mult1/result[4]~FF .SR_VALUE = 1'b0;
    defparam \mult1/result[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/result[5]~FF  (.D(\mult1/mult1/n127 ), .CE(ceg_net913), 
           .CLK(\clk~O ), .SR(resetn), .Q(\mult1/result[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/result[5]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/result[5]~FF .CE_POLARITY = 1'b0;
    defparam \mult1/result[5]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/result[5]~FF .D_POLARITY = 1'b1;
    defparam \mult1/result[5]~FF .SR_SYNC = 1'b0;
    defparam \mult1/result[5]~FF .SR_VALUE = 1'b0;
    defparam \mult1/result[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/result[6]~FF  (.D(\mult1/mult1/n126 ), .CE(ceg_net913), 
           .CLK(\clk~O ), .SR(resetn), .Q(\mult1/result[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/result[6]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/result[6]~FF .CE_POLARITY = 1'b0;
    defparam \mult1/result[6]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/result[6]~FF .D_POLARITY = 1'b1;
    defparam \mult1/result[6]~FF .SR_SYNC = 1'b0;
    defparam \mult1/result[6]~FF .SR_VALUE = 1'b0;
    defparam \mult1/result[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/result[7]~FF  (.D(\mult1/mult1/n125 ), .CE(ceg_net913), 
           .CLK(\clk~O ), .SR(resetn), .Q(\mult1/result[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/result[7]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/result[7]~FF .CE_POLARITY = 1'b0;
    defparam \mult1/result[7]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/result[7]~FF .D_POLARITY = 1'b1;
    defparam \mult1/result[7]~FF .SR_SYNC = 1'b0;
    defparam \mult1/result[7]~FF .SR_VALUE = 1'b0;
    defparam \mult1/result[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/result[8]~FF  (.D(\mult1/mult1/n124 ), .CE(ceg_net913), 
           .CLK(\clk~O ), .SR(resetn), .Q(\mult1/result[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/result[8]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/result[8]~FF .CE_POLARITY = 1'b0;
    defparam \mult1/result[8]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/result[8]~FF .D_POLARITY = 1'b1;
    defparam \mult1/result[8]~FF .SR_SYNC = 1'b0;
    defparam \mult1/result[8]~FF .SR_VALUE = 1'b0;
    defparam \mult1/result[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/result[9]~FF  (.D(\mult1/mult1/n123 ), .CE(ceg_net913), 
           .CLK(\clk~O ), .SR(resetn), .Q(\mult1/result[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/result[9]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/result[9]~FF .CE_POLARITY = 1'b0;
    defparam \mult1/result[9]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/result[9]~FF .D_POLARITY = 1'b1;
    defparam \mult1/result[9]~FF .SR_SYNC = 1'b0;
    defparam \mult1/result[9]~FF .SR_VALUE = 1'b0;
    defparam \mult1/result[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/result[10]~FF  (.D(\mult1/mult1/n122 ), .CE(ceg_net913), 
           .CLK(\clk~O ), .SR(resetn), .Q(\mult1/result[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/result[10]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/result[10]~FF .CE_POLARITY = 1'b0;
    defparam \mult1/result[10]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/result[10]~FF .D_POLARITY = 1'b1;
    defparam \mult1/result[10]~FF .SR_SYNC = 1'b0;
    defparam \mult1/result[10]~FF .SR_VALUE = 1'b0;
    defparam \mult1/result[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/result[11]~FF  (.D(\mult1/mult1/n121 ), .CE(ceg_net913), 
           .CLK(\clk~O ), .SR(resetn), .Q(\mult1/result[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/result[11]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/result[11]~FF .CE_POLARITY = 1'b0;
    defparam \mult1/result[11]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/result[11]~FF .D_POLARITY = 1'b1;
    defparam \mult1/result[11]~FF .SR_SYNC = 1'b0;
    defparam \mult1/result[11]~FF .SR_VALUE = 1'b0;
    defparam \mult1/result[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/result[12]~FF  (.D(\mult1/mult1/n120 ), .CE(ceg_net913), 
           .CLK(\clk~O ), .SR(resetn), .Q(\mult1/result[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/result[12]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/result[12]~FF .CE_POLARITY = 1'b0;
    defparam \mult1/result[12]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/result[12]~FF .D_POLARITY = 1'b1;
    defparam \mult1/result[12]~FF .SR_SYNC = 1'b0;
    defparam \mult1/result[12]~FF .SR_VALUE = 1'b0;
    defparam \mult1/result[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/result[13]~FF  (.D(\mult1/mult1/n119 ), .CE(ceg_net913), 
           .CLK(\clk~O ), .SR(resetn), .Q(\mult1/result[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/result[13]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/result[13]~FF .CE_POLARITY = 1'b0;
    defparam \mult1/result[13]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/result[13]~FF .D_POLARITY = 1'b1;
    defparam \mult1/result[13]~FF .SR_SYNC = 1'b0;
    defparam \mult1/result[13]~FF .SR_VALUE = 1'b0;
    defparam \mult1/result[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/result[14]~FF  (.D(\mult1/mult1/n118 ), .CE(ceg_net913), 
           .CLK(\clk~O ), .SR(resetn), .Q(\mult1/result[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/result[14]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/result[14]~FF .CE_POLARITY = 1'b0;
    defparam \mult1/result[14]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/result[14]~FF .D_POLARITY = 1'b1;
    defparam \mult1/result[14]~FF .SR_SYNC = 1'b0;
    defparam \mult1/result[14]~FF .SR_VALUE = 1'b0;
    defparam \mult1/result[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/result[15]~FF  (.D(\mult1/mult1/n117 ), .CE(ceg_net913), 
           .CLK(\clk~O ), .SR(resetn), .Q(\mult1/result[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/result[15]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/result[15]~FF .CE_POLARITY = 1'b0;
    defparam \mult1/result[15]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/result[15]~FF .D_POLARITY = 1'b1;
    defparam \mult1/result[15]~FF .SR_SYNC = 1'b0;
    defparam \mult1/result[15]~FF .SR_VALUE = 1'b0;
    defparam \mult1/result[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/result[16]~FF  (.D(\mult1/mult1/n116 ), .CE(ceg_net913), 
           .CLK(\clk~O ), .SR(resetn), .Q(\mult1/result[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/result[16]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/result[16]~FF .CE_POLARITY = 1'b0;
    defparam \mult1/result[16]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/result[16]~FF .D_POLARITY = 1'b1;
    defparam \mult1/result[16]~FF .SR_SYNC = 1'b0;
    defparam \mult1/result[16]~FF .SR_VALUE = 1'b0;
    defparam \mult1/result[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/result[17]~FF  (.D(\mult1/mult1/n115 ), .CE(ceg_net913), 
           .CLK(\clk~O ), .SR(resetn), .Q(\mult1/result[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/result[17]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/result[17]~FF .CE_POLARITY = 1'b0;
    defparam \mult1/result[17]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/result[17]~FF .D_POLARITY = 1'b1;
    defparam \mult1/result[17]~FF .SR_SYNC = 1'b0;
    defparam \mult1/result[17]~FF .SR_VALUE = 1'b0;
    defparam \mult1/result[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/result[18]~FF  (.D(\mult1/mult1/n114 ), .CE(ceg_net913), 
           .CLK(\clk~O ), .SR(resetn), .Q(\mult1/result[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/result[18]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/result[18]~FF .CE_POLARITY = 1'b0;
    defparam \mult1/result[18]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/result[18]~FF .D_POLARITY = 1'b1;
    defparam \mult1/result[18]~FF .SR_SYNC = 1'b0;
    defparam \mult1/result[18]~FF .SR_VALUE = 1'b0;
    defparam \mult1/result[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/result[19]~FF  (.D(\mult1/mult1/n113 ), .CE(ceg_net913), 
           .CLK(\clk~O ), .SR(resetn), .Q(\mult1/result[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/result[19]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/result[19]~FF .CE_POLARITY = 1'b0;
    defparam \mult1/result[19]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/result[19]~FF .D_POLARITY = 1'b1;
    defparam \mult1/result[19]~FF .SR_SYNC = 1'b0;
    defparam \mult1/result[19]~FF .SR_VALUE = 1'b0;
    defparam \mult1/result[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/result[20]~FF  (.D(\mult1/mult1/n112 ), .CE(ceg_net913), 
           .CLK(\clk~O ), .SR(resetn), .Q(\mult1/result[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/result[20]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/result[20]~FF .CE_POLARITY = 1'b0;
    defparam \mult1/result[20]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/result[20]~FF .D_POLARITY = 1'b1;
    defparam \mult1/result[20]~FF .SR_SYNC = 1'b0;
    defparam \mult1/result[20]~FF .SR_VALUE = 1'b0;
    defparam \mult1/result[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/result[21]~FF  (.D(\mult1/mult1/n111 ), .CE(ceg_net913), 
           .CLK(\clk~O ), .SR(resetn), .Q(\mult1/result[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/result[21]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/result[21]~FF .CE_POLARITY = 1'b0;
    defparam \mult1/result[21]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/result[21]~FF .D_POLARITY = 1'b1;
    defparam \mult1/result[21]~FF .SR_SYNC = 1'b0;
    defparam \mult1/result[21]~FF .SR_VALUE = 1'b0;
    defparam \mult1/result[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/result[22]~FF  (.D(\mult1/mult1/n110 ), .CE(ceg_net913), 
           .CLK(\clk~O ), .SR(resetn), .Q(\mult1/result[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/result[22]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/result[22]~FF .CE_POLARITY = 1'b0;
    defparam \mult1/result[22]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/result[22]~FF .D_POLARITY = 1'b1;
    defparam \mult1/result[22]~FF .SR_SYNC = 1'b0;
    defparam \mult1/result[22]~FF .SR_VALUE = 1'b0;
    defparam \mult1/result[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/result[23]~FF  (.D(\mult1/mult1/n109 ), .CE(ceg_net913), 
           .CLK(\clk~O ), .SR(resetn), .Q(\mult1/result[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/result[23]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/result[23]~FF .CE_POLARITY = 1'b0;
    defparam \mult1/result[23]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/result[23]~FF .D_POLARITY = 1'b1;
    defparam \mult1/result[23]~FF .SR_SYNC = 1'b0;
    defparam \mult1/result[23]~FF .SR_VALUE = 1'b0;
    defparam \mult1/result[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/result[24]~FF  (.D(\mult1/mult1/n108 ), .CE(ceg_net913), 
           .CLK(\clk~O ), .SR(resetn), .Q(\mult1/result[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/result[24]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/result[24]~FF .CE_POLARITY = 1'b0;
    defparam \mult1/result[24]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/result[24]~FF .D_POLARITY = 1'b1;
    defparam \mult1/result[24]~FF .SR_SYNC = 1'b0;
    defparam \mult1/result[24]~FF .SR_VALUE = 1'b0;
    defparam \mult1/result[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/result[25]~FF  (.D(\mult1/mult1/n107 ), .CE(ceg_net913), 
           .CLK(\clk~O ), .SR(resetn), .Q(\mult1/result[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/result[25]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/result[25]~FF .CE_POLARITY = 1'b0;
    defparam \mult1/result[25]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/result[25]~FF .D_POLARITY = 1'b1;
    defparam \mult1/result[25]~FF .SR_SYNC = 1'b0;
    defparam \mult1/result[25]~FF .SR_VALUE = 1'b0;
    defparam \mult1/result[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/result[26]~FF  (.D(\mult1/mult1/n106 ), .CE(ceg_net913), 
           .CLK(\clk~O ), .SR(resetn), .Q(\mult1/result[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/result[26]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/result[26]~FF .CE_POLARITY = 1'b0;
    defparam \mult1/result[26]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/result[26]~FF .D_POLARITY = 1'b1;
    defparam \mult1/result[26]~FF .SR_SYNC = 1'b0;
    defparam \mult1/result[26]~FF .SR_VALUE = 1'b0;
    defparam \mult1/result[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/result[27]~FF  (.D(\mult1/mult1/n105 ), .CE(ceg_net913), 
           .CLK(\clk~O ), .SR(resetn), .Q(\mult1/result[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/result[27]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/result[27]~FF .CE_POLARITY = 1'b0;
    defparam \mult1/result[27]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/result[27]~FF .D_POLARITY = 1'b1;
    defparam \mult1/result[27]~FF .SR_SYNC = 1'b0;
    defparam \mult1/result[27]~FF .SR_VALUE = 1'b0;
    defparam \mult1/result[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/result[28]~FF  (.D(\mult1/mult1/n104 ), .CE(ceg_net913), 
           .CLK(\clk~O ), .SR(resetn), .Q(\mult1/result[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/result[28]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/result[28]~FF .CE_POLARITY = 1'b0;
    defparam \mult1/result[28]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/result[28]~FF .D_POLARITY = 1'b1;
    defparam \mult1/result[28]~FF .SR_SYNC = 1'b0;
    defparam \mult1/result[28]~FF .SR_VALUE = 1'b0;
    defparam \mult1/result[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/result[29]~FF  (.D(\mult1/mult1/n103 ), .CE(ceg_net913), 
           .CLK(\clk~O ), .SR(resetn), .Q(\mult1/result[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/result[29]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/result[29]~FF .CE_POLARITY = 1'b0;
    defparam \mult1/result[29]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/result[29]~FF .D_POLARITY = 1'b1;
    defparam \mult1/result[29]~FF .SR_SYNC = 1'b0;
    defparam \mult1/result[29]~FF .SR_VALUE = 1'b0;
    defparam \mult1/result[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/result[30]~FF  (.D(\mult1/mult1/n102 ), .CE(ceg_net913), 
           .CLK(\clk~O ), .SR(resetn), .Q(\mult1/result[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/result[30]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/result[30]~FF .CE_POLARITY = 1'b0;
    defparam \mult1/result[30]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/result[30]~FF .D_POLARITY = 1'b1;
    defparam \mult1/result[30]~FF .SR_SYNC = 1'b0;
    defparam \mult1/result[30]~FF .SR_VALUE = 1'b0;
    defparam \mult1/result[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/result[31]~FF  (.D(\mult1/mult1/n101 ), .CE(ceg_net913), 
           .CLK(\clk~O ), .SR(resetn), .Q(\mult1/result[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/result[31]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/result[31]~FF .CE_POLARITY = 1'b0;
    defparam \mult1/result[31]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/result[31]~FF .D_POLARITY = 1'b1;
    defparam \mult1/result[31]~FF .SR_SYNC = 1'b0;
    defparam \mult1/result[31]~FF .SR_VALUE = 1'b0;
    defparam \mult1/result[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/state[1]~FF  (.D(\mult1/mult1/n63 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(resetn), .Q(\mult1/mult1/state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/state[1]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/state[1]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/mult1/state[1]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/state[1]~FF .SR_SYNC = 1'b0;
    defparam \mult1/mult1/state[1]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/state[2]~FF  (.D(\mult1/mult1/n62 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(resetn), .Q(\mult1/mult1/state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/state[2]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/state[2]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/state[2]~FF .SR_POLARITY = 1'b0;
    defparam \mult1/mult1/state[2]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/state[2]~FF .SR_SYNC = 1'b0;
    defparam \mult1/mult1/state[2]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/state[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/A[1]~FF  (.D(\mult1/mult1/n80 ), .CE(ceg_net839), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/A[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/A[1]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/A[1]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/A[1]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/A[1]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/A[1]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/A[1]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/A[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/A[2]~FF  (.D(\mult1/mult1/n79 ), .CE(ceg_net839), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/A[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/A[2]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/A[2]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/A[2]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/A[2]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/A[2]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/A[2]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/A[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/A[3]~FF  (.D(\mult1/mult1/n78 ), .CE(ceg_net839), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/A[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/A[3]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/A[3]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/A[3]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/A[3]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/A[3]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/A[3]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/A[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/A[4]~FF  (.D(\mult1/mult1/n77 ), .CE(ceg_net839), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/A[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/A[4]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/A[4]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/A[4]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/A[4]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/A[4]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/A[4]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/A[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/A[5]~FF  (.D(\mult1/mult1/n76 ), .CE(ceg_net839), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/A[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/A[5]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/A[5]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/A[5]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/A[5]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/A[5]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/A[5]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/A[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/A[6]~FF  (.D(\mult1/mult1/n75 ), .CE(ceg_net839), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/A[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/A[6]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/A[6]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/A[6]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/A[6]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/A[6]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/A[6]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/A[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/A[7]~FF  (.D(\mult1/mult1/n74 ), .CE(ceg_net839), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/A[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/A[7]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/A[7]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/A[7]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/A[7]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/A[7]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/A[7]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/A[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/A[8]~FF  (.D(\mult1/mult1/n73 ), .CE(ceg_net839), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/A[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/A[8]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/A[8]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/A[8]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/A[8]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/A[8]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/A[8]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/A[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/A[9]~FF  (.D(\mult1/mult1/n72 ), .CE(ceg_net839), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/A[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/A[9]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/A[9]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/A[9]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/A[9]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/A[9]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/A[9]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/A[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/A[10]~FF  (.D(\mult1/mult1/n71 ), .CE(ceg_net839), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/A[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/A[10]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/A[10]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/A[10]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/A[10]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/A[10]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/A[10]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/A[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/A[11]~FF  (.D(\mult1/mult1/n70 ), .CE(ceg_net839), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/A[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/A[11]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/A[11]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/A[11]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/A[11]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/A[11]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/A[11]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/A[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/A[12]~FF  (.D(\mult1/mult1/n69 ), .CE(ceg_net839), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/A[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/A[12]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/A[12]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/A[12]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/A[12]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/A[12]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/A[12]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/A[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/A[13]~FF  (.D(\mult1/mult1/n68 ), .CE(ceg_net839), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/A[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/A[13]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/A[13]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/A[13]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/A[13]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/A[13]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/A[13]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/A[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/A[14]~FF  (.D(\mult1/mult1/n67 ), .CE(ceg_net839), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/A[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/A[14]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/A[14]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/A[14]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/A[14]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/A[14]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/A[14]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/A[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/A[15]~FF  (.D(\mult1/mult1/n66 ), .CE(ceg_net839), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/A[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/A[15]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/A[15]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/A[15]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/A[15]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/A[15]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/A[15]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/A[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/B[1]~FF  (.D(\mult1/mult1/n97 ), .CE(ceg_net839), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/B[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/B[1]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/B[1]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/B[1]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/B[1]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/B[1]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/B[1]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/B[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/B[2]~FF  (.D(\mult1/mult1/n96 ), .CE(ceg_net839), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/B[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/B[2]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/B[2]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/B[2]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/B[2]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/B[2]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/B[2]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/B[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/B[3]~FF  (.D(\mult1/mult1/n95 ), .CE(ceg_net839), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/B[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/B[3]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/B[3]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/B[3]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/B[3]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/B[3]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/B[3]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/B[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/B[4]~FF  (.D(\mult1/mult1/n94 ), .CE(ceg_net839), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/B[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/B[4]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/B[4]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/B[4]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/B[4]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/B[4]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/B[4]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/B[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/B[5]~FF  (.D(\mult1/mult1/n93 ), .CE(ceg_net839), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/B[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/B[5]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/B[5]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/B[5]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/B[5]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/B[5]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/B[5]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/B[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/B[6]~FF  (.D(\mult1/mult1/n92 ), .CE(ceg_net839), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/B[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/B[6]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/B[6]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/B[6]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/B[6]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/B[6]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/B[6]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/B[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/B[7]~FF  (.D(\mult1/mult1/n91 ), .CE(ceg_net839), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/B[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/B[7]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/B[7]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/B[7]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/B[7]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/B[7]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/B[7]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/B[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/B[8]~FF  (.D(\mult1/mult1/n90 ), .CE(ceg_net839), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/B[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/B[8]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/B[8]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/B[8]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/B[8]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/B[8]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/B[8]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/B[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/B[9]~FF  (.D(\mult1/mult1/n89 ), .CE(ceg_net839), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/B[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/B[9]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/B[9]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/B[9]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/B[9]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/B[9]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/B[9]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/B[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/B[10]~FF  (.D(\mult1/mult1/n88 ), .CE(ceg_net839), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/B[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/B[10]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/B[10]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/B[10]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/B[10]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/B[10]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/B[10]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/B[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/B[11]~FF  (.D(\mult1/mult1/n87 ), .CE(ceg_net839), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/B[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/B[11]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/B[11]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/B[11]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/B[11]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/B[11]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/B[11]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/B[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/B[12]~FF  (.D(\mult1/mult1/n86 ), .CE(ceg_net839), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/B[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/B[12]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/B[12]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/B[12]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/B[12]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/B[12]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/B[12]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/B[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/B[13]~FF  (.D(\mult1/mult1/n85 ), .CE(ceg_net839), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/B[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/B[13]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/B[13]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/B[13]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/B[13]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/B[13]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/B[13]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/B[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/B[14]~FF  (.D(\mult1/mult1/n84 ), .CE(ceg_net839), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/B[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/B[14]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/B[14]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/B[14]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/B[14]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/B[14]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/B[14]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/B[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/B[15]~FF  (.D(\mult1/mult1/n83 ), .CE(ceg_net839), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/B[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/B[15]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/B[15]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/B[15]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/B[15]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/B[15]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/B[15]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/B[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/count[1]~FF  (.D(\mult1/mult1/n137 ), .CE(ceg_net847), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/count[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/count[1]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/count[1]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/count[1]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/count[1]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/count[1]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/count[1]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/count[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/count[2]~FF  (.D(\mult1/mult1/n136 ), .CE(ceg_net847), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/count[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/count[2]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/count[2]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/count[2]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/count[2]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/count[2]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/count[2]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/count[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/count[3]~FF  (.D(\mult1/mult1/n135 ), .CE(ceg_net847), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/count[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/count[3]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/count[3]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/count[3]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/count[3]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/count[3]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/count[3]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/count[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \mult1/mult1/count[4]~FF  (.D(\mult1/mult1/n134 ), .CE(ceg_net847), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\mult1/mult1/count[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(90)
    defparam \mult1/mult1/count[4]~FF .CLK_POLARITY = 1'b1;
    defparam \mult1/mult1/count[4]~FF .CE_POLARITY = 1'b1;
    defparam \mult1/mult1/count[4]~FF .SR_POLARITY = 1'b1;
    defparam \mult1/mult1/count[4]~FF .D_POLARITY = 1'b1;
    defparam \mult1/mult1/count[4]~FF .SR_SYNC = 1'b1;
    defparam \mult1/mult1/count[4]~FF .SR_VALUE = 1'b0;
    defparam \mult1/mult1/count[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_ADD \CPU/add_33/i1  (.I0(n1587), .I1(\CPU/rs1[0] ), .CI(1'b0), 
            .O(n6), .CO(n7)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(131)
    defparam \CPU/add_33/i1 .I0_POLARITY = 1'b0;
    defparam \CPU/add_33/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_90/i2  (.I0(\CPU/PC[1] ), .I1(n787), .CI(1'b0), .O(n8), 
            .CO(n9)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(207)
    defparam \CPU/add_90/i2 .I0_POLARITY = 1'b1;
    defparam \CPU/add_90/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_92/i1  (.I0(\CPU/rs1[0] ), .I1(n793), .CI(1'b0), 
            .O(n12), .CO(n13)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(212)
    defparam \CPU/add_92/i1 .I0_POLARITY = 1'b1;
    defparam \CPU/add_92/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_603/i1  (.I0(\CPU/cycles[1] ), .I1(\CPU/cycles[0] ), 
            .CI(1'b0), .O(n14), .CO(n15)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/add_603/i1 .I0_POLARITY = 1'b1;
    defparam \CPU/add_603/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \mult1/mult1/add_8/i1  (.I0(\mult1/result[0] ), .I1(\mult1/mult1/A[0] ), 
            .CI(1'b0), .O(n209), .CO(n210)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(76)
    defparam \mult1/mult1/add_8/i1 .I0_POLARITY = 1'b1;
    defparam \mult1/mult1/add_8/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \mult1/mult1/add_8/i2  (.I0(\mult1/result[1] ), .I1(\mult1/mult1/A[1] ), 
            .CI(n210), .O(n238), .CO(n239)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(76)
    defparam \mult1/mult1/add_8/i2 .I0_POLARITY = 1'b1;
    defparam \mult1/mult1/add_8/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \mult1/mult1/add_8/i32  (.I0(\mult1/result[31] ), .I1(1'b0), 
            .CI(n453), .O(n451)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(76)
    defparam \mult1/mult1/add_8/i32 .I0_POLARITY = 1'b1;
    defparam \mult1/mult1/add_8/i32 .I1_POLARITY = 1'b1;
    EFX_ADD \mult1/mult1/add_8/i31  (.I0(\mult1/result[30] ), .I1(1'b0), 
            .CI(n455), .O(n452), .CO(n453)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(76)
    defparam \mult1/mult1/add_8/i31 .I0_POLARITY = 1'b1;
    defparam \mult1/mult1/add_8/i31 .I1_POLARITY = 1'b1;
    EFX_ADD \mult1/mult1/add_8/i30  (.I0(\mult1/result[29] ), .I1(1'b0), 
            .CI(n457), .O(n454), .CO(n455)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(76)
    defparam \mult1/mult1/add_8/i30 .I0_POLARITY = 1'b1;
    defparam \mult1/mult1/add_8/i30 .I1_POLARITY = 1'b1;
    EFX_ADD \mult1/mult1/add_8/i29  (.I0(\mult1/result[28] ), .I1(1'b0), 
            .CI(n459), .O(n456), .CO(n457)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(76)
    defparam \mult1/mult1/add_8/i29 .I0_POLARITY = 1'b1;
    defparam \mult1/mult1/add_8/i29 .I1_POLARITY = 1'b1;
    EFX_ADD \mult1/mult1/add_8/i28  (.I0(\mult1/result[27] ), .I1(1'b0), 
            .CI(n461), .O(n458), .CO(n459)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(76)
    defparam \mult1/mult1/add_8/i28 .I0_POLARITY = 1'b1;
    defparam \mult1/mult1/add_8/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \mult1/mult1/add_8/i27  (.I0(\mult1/result[26] ), .I1(1'b0), 
            .CI(n463), .O(n460), .CO(n461)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(76)
    defparam \mult1/mult1/add_8/i27 .I0_POLARITY = 1'b1;
    defparam \mult1/mult1/add_8/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \mult1/mult1/add_8/i26  (.I0(\mult1/result[25] ), .I1(1'b0), 
            .CI(n465), .O(n462), .CO(n463)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(76)
    defparam \mult1/mult1/add_8/i26 .I0_POLARITY = 1'b1;
    defparam \mult1/mult1/add_8/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \mult1/mult1/add_8/i25  (.I0(\mult1/result[24] ), .I1(1'b0), 
            .CI(n467), .O(n464), .CO(n465)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(76)
    defparam \mult1/mult1/add_8/i25 .I0_POLARITY = 1'b1;
    defparam \mult1/mult1/add_8/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \mult1/mult1/add_8/i24  (.I0(\mult1/result[23] ), .I1(1'b0), 
            .CI(n469), .O(n466), .CO(n467)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(76)
    defparam \mult1/mult1/add_8/i24 .I0_POLARITY = 1'b1;
    defparam \mult1/mult1/add_8/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \mult1/mult1/add_8/i23  (.I0(\mult1/result[22] ), .I1(1'b0), 
            .CI(n471), .O(n468), .CO(n469)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(76)
    defparam \mult1/mult1/add_8/i23 .I0_POLARITY = 1'b1;
    defparam \mult1/mult1/add_8/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \mult1/mult1/add_8/i22  (.I0(\mult1/result[21] ), .I1(1'b0), 
            .CI(n473), .O(n470), .CO(n471)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(76)
    defparam \mult1/mult1/add_8/i22 .I0_POLARITY = 1'b1;
    defparam \mult1/mult1/add_8/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \mult1/mult1/add_8/i21  (.I0(\mult1/result[20] ), .I1(1'b0), 
            .CI(n475), .O(n472), .CO(n473)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(76)
    defparam \mult1/mult1/add_8/i21 .I0_POLARITY = 1'b1;
    defparam \mult1/mult1/add_8/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \mult1/mult1/add_8/i20  (.I0(\mult1/result[19] ), .I1(1'b0), 
            .CI(n477), .O(n474), .CO(n475)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(76)
    defparam \mult1/mult1/add_8/i20 .I0_POLARITY = 1'b1;
    defparam \mult1/mult1/add_8/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \mult1/mult1/add_8/i19  (.I0(\mult1/result[18] ), .I1(1'b0), 
            .CI(n479), .O(n476), .CO(n477)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(76)
    defparam \mult1/mult1/add_8/i19 .I0_POLARITY = 1'b1;
    defparam \mult1/mult1/add_8/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \mult1/mult1/add_8/i18  (.I0(\mult1/result[17] ), .I1(1'b0), 
            .CI(n481), .O(n478), .CO(n479)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(76)
    defparam \mult1/mult1/add_8/i18 .I0_POLARITY = 1'b1;
    defparam \mult1/mult1/add_8/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \mult1/mult1/add_8/i17  (.I0(\mult1/result[16] ), .I1(1'b0), 
            .CI(n483), .O(n480), .CO(n481)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(76)
    defparam \mult1/mult1/add_8/i17 .I0_POLARITY = 1'b1;
    defparam \mult1/mult1/add_8/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \mult1/mult1/add_8/i16  (.I0(\mult1/result[15] ), .I1(\mult1/mult1/A[15] ), 
            .CI(n485), .O(n482), .CO(n483)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(76)
    defparam \mult1/mult1/add_8/i16 .I0_POLARITY = 1'b1;
    defparam \mult1/mult1/add_8/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \mult1/mult1/add_8/i15  (.I0(\mult1/result[14] ), .I1(\mult1/mult1/A[14] ), 
            .CI(n487), .O(n484), .CO(n485)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(76)
    defparam \mult1/mult1/add_8/i15 .I0_POLARITY = 1'b1;
    defparam \mult1/mult1/add_8/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \mult1/mult1/add_8/i14  (.I0(\mult1/result[13] ), .I1(\mult1/mult1/A[13] ), 
            .CI(n489), .O(n486), .CO(n487)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(76)
    defparam \mult1/mult1/add_8/i14 .I0_POLARITY = 1'b1;
    defparam \mult1/mult1/add_8/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \mult1/mult1/add_8/i13  (.I0(\mult1/result[12] ), .I1(\mult1/mult1/A[12] ), 
            .CI(n491), .O(n488), .CO(n489)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(76)
    defparam \mult1/mult1/add_8/i13 .I0_POLARITY = 1'b1;
    defparam \mult1/mult1/add_8/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \mult1/mult1/add_8/i12  (.I0(\mult1/result[11] ), .I1(\mult1/mult1/A[11] ), 
            .CI(n493), .O(n490), .CO(n491)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(76)
    defparam \mult1/mult1/add_8/i12 .I0_POLARITY = 1'b1;
    defparam \mult1/mult1/add_8/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \mult1/mult1/add_8/i11  (.I0(\mult1/result[10] ), .I1(\mult1/mult1/A[10] ), 
            .CI(n495), .O(n492), .CO(n493)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(76)
    defparam \mult1/mult1/add_8/i11 .I0_POLARITY = 1'b1;
    defparam \mult1/mult1/add_8/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \mult1/mult1/add_8/i10  (.I0(\mult1/result[9] ), .I1(\mult1/mult1/A[9] ), 
            .CI(n497), .O(n494), .CO(n495)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(76)
    defparam \mult1/mult1/add_8/i10 .I0_POLARITY = 1'b1;
    defparam \mult1/mult1/add_8/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \mult1/mult1/add_8/i9  (.I0(\mult1/result[8] ), .I1(\mult1/mult1/A[8] ), 
            .CI(n499), .O(n496), .CO(n497)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(76)
    defparam \mult1/mult1/add_8/i9 .I0_POLARITY = 1'b1;
    defparam \mult1/mult1/add_8/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \mult1/mult1/add_8/i8  (.I0(\mult1/result[7] ), .I1(\mult1/mult1/A[7] ), 
            .CI(n501), .O(n498), .CO(n499)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(76)
    defparam \mult1/mult1/add_8/i8 .I0_POLARITY = 1'b1;
    defparam \mult1/mult1/add_8/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \mult1/mult1/add_8/i7  (.I0(\mult1/result[6] ), .I1(\mult1/mult1/A[6] ), 
            .CI(n503), .O(n500), .CO(n501)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(76)
    defparam \mult1/mult1/add_8/i7 .I0_POLARITY = 1'b1;
    defparam \mult1/mult1/add_8/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \mult1/mult1/add_8/i6  (.I0(\mult1/result[5] ), .I1(\mult1/mult1/A[5] ), 
            .CI(n505), .O(n502), .CO(n503)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(76)
    defparam \mult1/mult1/add_8/i6 .I0_POLARITY = 1'b1;
    defparam \mult1/mult1/add_8/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \mult1/mult1/add_8/i5  (.I0(\mult1/result[4] ), .I1(\mult1/mult1/A[4] ), 
            .CI(n507), .O(n504), .CO(n505)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(76)
    defparam \mult1/mult1/add_8/i5 .I0_POLARITY = 1'b1;
    defparam \mult1/mult1/add_8/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \mult1/mult1/add_8/i4  (.I0(\mult1/result[3] ), .I1(\mult1/mult1/A[3] ), 
            .CI(n509), .O(n506), .CO(n507)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(76)
    defparam \mult1/mult1/add_8/i4 .I0_POLARITY = 1'b1;
    defparam \mult1/mult1/add_8/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \mult1/mult1/add_8/i3  (.I0(\mult1/result[2] ), .I1(\mult1/mult1/A[2] ), 
            .CI(n239), .O(n508), .CO(n509)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/mult/mult.v(76)
    defparam \mult1/mult1/add_8/i3 .I0_POLARITY = 1'b1;
    defparam \mult1/mult1/add_8/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_603/i31  (.I0(\CPU/cycles[31] ), .I1(1'b0), .CI(n512), 
            .O(n510)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/add_603/i31 .I0_POLARITY = 1'b1;
    defparam \CPU/add_603/i31 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_603/i30  (.I0(\CPU/cycles[30] ), .I1(1'b0), .CI(n514), 
            .O(n511), .CO(n512)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/add_603/i30 .I0_POLARITY = 1'b1;
    defparam \CPU/add_603/i30 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_603/i29  (.I0(\CPU/cycles[29] ), .I1(1'b0), .CI(n516), 
            .O(n513), .CO(n514)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/add_603/i29 .I0_POLARITY = 1'b1;
    defparam \CPU/add_603/i29 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_603/i28  (.I0(\CPU/cycles[28] ), .I1(1'b0), .CI(n518), 
            .O(n515), .CO(n516)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/add_603/i28 .I0_POLARITY = 1'b1;
    defparam \CPU/add_603/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_603/i27  (.I0(\CPU/cycles[27] ), .I1(1'b0), .CI(n520), 
            .O(n517), .CO(n518)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/add_603/i27 .I0_POLARITY = 1'b1;
    defparam \CPU/add_603/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_603/i26  (.I0(\CPU/cycles[26] ), .I1(1'b0), .CI(n522), 
            .O(n519), .CO(n520)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/add_603/i26 .I0_POLARITY = 1'b1;
    defparam \CPU/add_603/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_603/i25  (.I0(\CPU/cycles[25] ), .I1(1'b0), .CI(n524), 
            .O(n521), .CO(n522)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/add_603/i25 .I0_POLARITY = 1'b1;
    defparam \CPU/add_603/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_603/i24  (.I0(\CPU/cycles[24] ), .I1(1'b0), .CI(n526), 
            .O(n523), .CO(n524)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/add_603/i24 .I0_POLARITY = 1'b1;
    defparam \CPU/add_603/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_603/i23  (.I0(\CPU/cycles[23] ), .I1(1'b0), .CI(n528), 
            .O(n525), .CO(n526)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/add_603/i23 .I0_POLARITY = 1'b1;
    defparam \CPU/add_603/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_603/i22  (.I0(\CPU/cycles[22] ), .I1(1'b0), .CI(n530), 
            .O(n527), .CO(n528)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/add_603/i22 .I0_POLARITY = 1'b1;
    defparam \CPU/add_603/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_603/i21  (.I0(\CPU/cycles[21] ), .I1(1'b0), .CI(n532), 
            .O(n529), .CO(n530)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/add_603/i21 .I0_POLARITY = 1'b1;
    defparam \CPU/add_603/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_603/i20  (.I0(\CPU/cycles[20] ), .I1(1'b0), .CI(n534), 
            .O(n531), .CO(n532)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/add_603/i20 .I0_POLARITY = 1'b1;
    defparam \CPU/add_603/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_603/i19  (.I0(\CPU/cycles[19] ), .I1(1'b0), .CI(n536), 
            .O(n533), .CO(n534)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/add_603/i19 .I0_POLARITY = 1'b1;
    defparam \CPU/add_603/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_603/i18  (.I0(\CPU/cycles[18] ), .I1(1'b0), .CI(n538), 
            .O(n535), .CO(n536)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/add_603/i18 .I0_POLARITY = 1'b1;
    defparam \CPU/add_603/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_603/i17  (.I0(\CPU/cycles[17] ), .I1(1'b0), .CI(n540), 
            .O(n537), .CO(n538)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/add_603/i17 .I0_POLARITY = 1'b1;
    defparam \CPU/add_603/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_603/i16  (.I0(\CPU/cycles[16] ), .I1(1'b0), .CI(n542), 
            .O(n539), .CO(n540)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/add_603/i16 .I0_POLARITY = 1'b1;
    defparam \CPU/add_603/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_603/i15  (.I0(\CPU/cycles[15] ), .I1(1'b0), .CI(n544), 
            .O(n541), .CO(n542)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/add_603/i15 .I0_POLARITY = 1'b1;
    defparam \CPU/add_603/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_603/i14  (.I0(\CPU/cycles[14] ), .I1(1'b0), .CI(n546), 
            .O(n543), .CO(n544)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/add_603/i14 .I0_POLARITY = 1'b1;
    defparam \CPU/add_603/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_603/i13  (.I0(\CPU/cycles[13] ), .I1(1'b0), .CI(n548), 
            .O(n545), .CO(n546)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/add_603/i13 .I0_POLARITY = 1'b1;
    defparam \CPU/add_603/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_603/i12  (.I0(\CPU/cycles[12] ), .I1(1'b0), .CI(n550), 
            .O(n547), .CO(n548)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/add_603/i12 .I0_POLARITY = 1'b1;
    defparam \CPU/add_603/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_603/i11  (.I0(\CPU/cycles[11] ), .I1(1'b0), .CI(n552), 
            .O(n549), .CO(n550)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/add_603/i11 .I0_POLARITY = 1'b1;
    defparam \CPU/add_603/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_603/i10  (.I0(\CPU/cycles[10] ), .I1(1'b0), .CI(n554), 
            .O(n551), .CO(n552)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/add_603/i10 .I0_POLARITY = 1'b1;
    defparam \CPU/add_603/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_603/i9  (.I0(\CPU/cycles[9] ), .I1(1'b0), .CI(n556), 
            .O(n553), .CO(n554)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/add_603/i9 .I0_POLARITY = 1'b1;
    defparam \CPU/add_603/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_603/i8  (.I0(\CPU/cycles[8] ), .I1(1'b0), .CI(n558), 
            .O(n555), .CO(n556)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/add_603/i8 .I0_POLARITY = 1'b1;
    defparam \CPU/add_603/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_603/i7  (.I0(\CPU/cycles[7] ), .I1(1'b0), .CI(n560), 
            .O(n557), .CO(n558)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/add_603/i7 .I0_POLARITY = 1'b1;
    defparam \CPU/add_603/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_603/i6  (.I0(\CPU/cycles[6] ), .I1(1'b0), .CI(n562), 
            .O(n559), .CO(n560)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/add_603/i6 .I0_POLARITY = 1'b1;
    defparam \CPU/add_603/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_603/i5  (.I0(\CPU/cycles[5] ), .I1(1'b0), .CI(n564), 
            .O(n561), .CO(n562)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/add_603/i5 .I0_POLARITY = 1'b1;
    defparam \CPU/add_603/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_603/i4  (.I0(\CPU/cycles[4] ), .I1(1'b0), .CI(n566), 
            .O(n563), .CO(n564)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/add_603/i4 .I0_POLARITY = 1'b1;
    defparam \CPU/add_603/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_603/i3  (.I0(\CPU/cycles[3] ), .I1(1'b0), .CI(n568), 
            .O(n565), .CO(n566)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/add_603/i3 .I0_POLARITY = 1'b1;
    defparam \CPU/add_603/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_603/i2  (.I0(\CPU/cycles[2] ), .I1(1'b0), .CI(n15), 
            .O(n567), .CO(n568)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(380)
    defparam \CPU/add_603/i2 .I0_POLARITY = 1'b1;
    defparam \CPU/add_603/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_92/i24  (.I0(\CPU/rs1[23] ), .I1(\CPU/instr[31] ), 
            .CI(n571), .O(n569)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(212)
    defparam \CPU/add_92/i24 .I0_POLARITY = 1'b1;
    defparam \CPU/add_92/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_92/i23  (.I0(\CPU/rs1[22] ), .I1(\CPU/instr[31] ), 
            .CI(n573), .O(n570), .CO(n571)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(212)
    defparam \CPU/add_92/i23 .I0_POLARITY = 1'b1;
    defparam \CPU/add_92/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_92/i22  (.I0(\CPU/rs1[21] ), .I1(\CPU/instr[31] ), 
            .CI(n575), .O(n572), .CO(n573)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(212)
    defparam \CPU/add_92/i22 .I0_POLARITY = 1'b1;
    defparam \CPU/add_92/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_92/i21  (.I0(\CPU/rs1[20] ), .I1(\CPU/instr[31] ), 
            .CI(n577), .O(n574), .CO(n575)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(212)
    defparam \CPU/add_92/i21 .I0_POLARITY = 1'b1;
    defparam \CPU/add_92/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_92/i20  (.I0(\CPU/rs1[19] ), .I1(\CPU/instr[31] ), 
            .CI(n579), .O(n576), .CO(n577)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(212)
    defparam \CPU/add_92/i20 .I0_POLARITY = 1'b1;
    defparam \CPU/add_92/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_92/i19  (.I0(\CPU/rs1[18] ), .I1(\CPU/instr[31] ), 
            .CI(n581), .O(n578), .CO(n579)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(212)
    defparam \CPU/add_92/i19 .I0_POLARITY = 1'b1;
    defparam \CPU/add_92/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_92/i18  (.I0(\CPU/rs1[17] ), .I1(\CPU/instr[31] ), 
            .CI(n583), .O(n580), .CO(n581)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(212)
    defparam \CPU/add_92/i18 .I0_POLARITY = 1'b1;
    defparam \CPU/add_92/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_92/i17  (.I0(\CPU/rs1[16] ), .I1(\CPU/instr[31] ), 
            .CI(n585), .O(n582), .CO(n583)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(212)
    defparam \CPU/add_92/i17 .I0_POLARITY = 1'b1;
    defparam \CPU/add_92/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_92/i16  (.I0(\CPU/rs1[15] ), .I1(\CPU/instr[31] ), 
            .CI(n587), .O(n584), .CO(n585)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(212)
    defparam \CPU/add_92/i16 .I0_POLARITY = 1'b1;
    defparam \CPU/add_92/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_92/i15  (.I0(\CPU/rs1[14] ), .I1(\CPU/instr[31] ), 
            .CI(n589), .O(n586), .CO(n587)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(212)
    defparam \CPU/add_92/i15 .I0_POLARITY = 1'b1;
    defparam \CPU/add_92/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_92/i14  (.I0(\CPU/rs1[13] ), .I1(\CPU/instr[31] ), 
            .CI(n591), .O(n588), .CO(n589)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(212)
    defparam \CPU/add_92/i14 .I0_POLARITY = 1'b1;
    defparam \CPU/add_92/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_92/i13  (.I0(\CPU/rs1[12] ), .I1(\CPU/instr[31] ), 
            .CI(n593), .O(n590), .CO(n591)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(212)
    defparam \CPU/add_92/i13 .I0_POLARITY = 1'b1;
    defparam \CPU/add_92/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_92/i12  (.I0(\CPU/rs1[11] ), .I1(\CPU/instr[31] ), 
            .CI(n595), .O(n592), .CO(n593)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(212)
    defparam \CPU/add_92/i12 .I0_POLARITY = 1'b1;
    defparam \CPU/add_92/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_92/i11  (.I0(\CPU/rs1[10] ), .I1(\CPU/instr[30] ), 
            .CI(n597), .O(n594), .CO(n595)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(212)
    defparam \CPU/add_92/i11 .I0_POLARITY = 1'b1;
    defparam \CPU/add_92/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_92/i10  (.I0(\CPU/rs1[9] ), .I1(\CPU/instr[29] ), .CI(n599), 
            .O(n596), .CO(n597)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(212)
    defparam \CPU/add_92/i10 .I0_POLARITY = 1'b1;
    defparam \CPU/add_92/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_92/i9  (.I0(\CPU/rs1[8] ), .I1(\CPU/instr[28] ), .CI(n601), 
            .O(n598), .CO(n599)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(212)
    defparam \CPU/add_92/i9 .I0_POLARITY = 1'b1;
    defparam \CPU/add_92/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_92/i8  (.I0(\CPU/rs1[7] ), .I1(\CPU/instr[27] ), .CI(n603), 
            .O(n600), .CO(n601)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(212)
    defparam \CPU/add_92/i8 .I0_POLARITY = 1'b1;
    defparam \CPU/add_92/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_92/i7  (.I0(\CPU/rs1[6] ), .I1(\CPU/instr[26] ), .CI(n605), 
            .O(n602), .CO(n603)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(212)
    defparam \CPU/add_92/i7 .I0_POLARITY = 1'b1;
    defparam \CPU/add_92/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_92/i6  (.I0(\CPU/rs1[5] ), .I1(\CPU/instr[25] ), .CI(n607), 
            .O(n604), .CO(n605)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(212)
    defparam \CPU/add_92/i6 .I0_POLARITY = 1'b1;
    defparam \CPU/add_92/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_92/i5  (.I0(\CPU/rs1[4] ), .I1(n1378), .CI(n609), 
            .O(n606), .CO(n607)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(212)
    defparam \CPU/add_92/i5 .I0_POLARITY = 1'b1;
    defparam \CPU/add_92/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_92/i4  (.I0(\CPU/rs1[3] ), .I1(n1381), .CI(n611), 
            .O(n608), .CO(n609)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(212)
    defparam \CPU/add_92/i4 .I0_POLARITY = 1'b1;
    defparam \CPU/add_92/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_92/i3  (.I0(\CPU/rs1[2] ), .I1(n1384), .CI(n613), 
            .O(n610), .CO(n611)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(212)
    defparam \CPU/add_92/i3 .I0_POLARITY = 1'b1;
    defparam \CPU/add_92/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_92/i2  (.I0(\CPU/rs1[1] ), .I1(n1387), .CI(n13), 
            .O(n612), .CO(n613)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(212)
    defparam \CPU/add_92/i2 .I0_POLARITY = 1'b1;
    defparam \CPU/add_92/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_90/i24  (.I0(\CPU/PC[23] ), .I1(n1390), .CI(n616), 
            .O(n614)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(207)
    defparam \CPU/add_90/i24 .I0_POLARITY = 1'b1;
    defparam \CPU/add_90/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_90/i23  (.I0(\CPU/PC[22] ), .I1(n1393), .CI(n618), 
            .O(n615), .CO(n616)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(207)
    defparam \CPU/add_90/i23 .I0_POLARITY = 1'b1;
    defparam \CPU/add_90/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_90/i22  (.I0(\CPU/PC[21] ), .I1(n1396), .CI(n620), 
            .O(n617), .CO(n618)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(207)
    defparam \CPU/add_90/i22 .I0_POLARITY = 1'b1;
    defparam \CPU/add_90/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_90/i21  (.I0(\CPU/PC[20] ), .I1(n1399), .CI(n622), 
            .O(n619), .CO(n620)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(207)
    defparam \CPU/add_90/i21 .I0_POLARITY = 1'b1;
    defparam \CPU/add_90/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_90/i20  (.I0(\CPU/PC[19] ), .I1(n1402), .CI(n624), 
            .O(n621), .CO(n622)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(207)
    defparam \CPU/add_90/i20 .I0_POLARITY = 1'b1;
    defparam \CPU/add_90/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_90/i19  (.I0(\CPU/PC[18] ), .I1(n1405), .CI(n626), 
            .O(n623), .CO(n624)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(207)
    defparam \CPU/add_90/i19 .I0_POLARITY = 1'b1;
    defparam \CPU/add_90/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_90/i18  (.I0(\CPU/PC[17] ), .I1(n1408), .CI(n628), 
            .O(n625), .CO(n626)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(207)
    defparam \CPU/add_90/i18 .I0_POLARITY = 1'b1;
    defparam \CPU/add_90/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_90/i17  (.I0(\CPU/PC[16] ), .I1(n1411), .CI(n630), 
            .O(n627), .CO(n628)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(207)
    defparam \CPU/add_90/i17 .I0_POLARITY = 1'b1;
    defparam \CPU/add_90/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_90/i16  (.I0(\CPU/PC[15] ), .I1(n1414), .CI(n632), 
            .O(n629), .CO(n630)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(207)
    defparam \CPU/add_90/i16 .I0_POLARITY = 1'b1;
    defparam \CPU/add_90/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_90/i15  (.I0(\CPU/PC[14] ), .I1(n1417), .CI(n634), 
            .O(n631), .CO(n632)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(207)
    defparam \CPU/add_90/i15 .I0_POLARITY = 1'b1;
    defparam \CPU/add_90/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_90/i14  (.I0(\CPU/PC[13] ), .I1(n1420), .CI(n636), 
            .O(n633), .CO(n634)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(207)
    defparam \CPU/add_90/i14 .I0_POLARITY = 1'b1;
    defparam \CPU/add_90/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_90/i13  (.I0(\CPU/PC[12] ), .I1(n1423), .CI(n638), 
            .O(n635), .CO(n636)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(207)
    defparam \CPU/add_90/i13 .I0_POLARITY = 1'b1;
    defparam \CPU/add_90/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_90/i12  (.I0(\CPU/PC[11] ), .I1(n1426), .CI(n640), 
            .O(n637), .CO(n638)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(207)
    defparam \CPU/add_90/i12 .I0_POLARITY = 1'b1;
    defparam \CPU/add_90/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_90/i11  (.I0(\CPU/PC[10] ), .I1(n1429), .CI(n642), 
            .O(n639), .CO(n640)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(207)
    defparam \CPU/add_90/i11 .I0_POLARITY = 1'b1;
    defparam \CPU/add_90/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_90/i10  (.I0(\CPU/PC[9] ), .I1(n1432), .CI(n644), 
            .O(n641), .CO(n642)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(207)
    defparam \CPU/add_90/i10 .I0_POLARITY = 1'b1;
    defparam \CPU/add_90/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_90/i9  (.I0(\CPU/PC[8] ), .I1(n1435), .CI(n646), 
            .O(n643), .CO(n644)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(207)
    defparam \CPU/add_90/i9 .I0_POLARITY = 1'b1;
    defparam \CPU/add_90/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_90/i8  (.I0(\CPU/PC[7] ), .I1(n1438), .CI(n648), 
            .O(n645), .CO(n646)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(207)
    defparam \CPU/add_90/i8 .I0_POLARITY = 1'b1;
    defparam \CPU/add_90/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_90/i7  (.I0(\CPU/PC[6] ), .I1(n1441), .CI(n650), 
            .O(n647), .CO(n648)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(207)
    defparam \CPU/add_90/i7 .I0_POLARITY = 1'b1;
    defparam \CPU/add_90/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_90/i6  (.I0(\CPU/PC[5] ), .I1(n1444), .CI(n652), 
            .O(n649), .CO(n650)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(207)
    defparam \CPU/add_90/i6 .I0_POLARITY = 1'b1;
    defparam \CPU/add_90/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_90/i5  (.I0(\CPU/PC[4] ), .I1(n1447), .CI(n654), 
            .O(n651), .CO(n652)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(207)
    defparam \CPU/add_90/i5 .I0_POLARITY = 1'b1;
    defparam \CPU/add_90/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_90/i4  (.I0(\CPU/PC[3] ), .I1(n1450), .CI(n656), 
            .O(n653), .CO(n654)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(207)
    defparam \CPU/add_90/i4 .I0_POLARITY = 1'b1;
    defparam \CPU/add_90/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_90/i3  (.I0(\CPU/PC[2] ), .I1(n1453), .CI(n9), .O(n655), 
            .CO(n656)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(207)
    defparam \CPU/add_90/i3 .I0_POLARITY = 1'b1;
    defparam \CPU/add_90/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_33/i32  (.I0(n1525), .I1(\CPU/rs1[31] ), .CI(n660), 
            .O(n657), .CO(n2159)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(131)
    defparam \CPU/add_33/i32 .I0_POLARITY = 1'b0;
    defparam \CPU/add_33/i32 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_33/i31  (.I0(n1527), .I1(\CPU/rs1[30] ), .CI(n662), 
            .O(n659), .CO(n660)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(131)
    defparam \CPU/add_33/i31 .I0_POLARITY = 1'b0;
    defparam \CPU/add_33/i31 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_33/i30  (.I0(n1529), .I1(\CPU/rs1[29] ), .CI(n664), 
            .O(n661), .CO(n662)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(131)
    defparam \CPU/add_33/i30 .I0_POLARITY = 1'b0;
    defparam \CPU/add_33/i30 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_33/i29  (.I0(n1531), .I1(\CPU/rs1[28] ), .CI(n666), 
            .O(n663), .CO(n664)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(131)
    defparam \CPU/add_33/i29 .I0_POLARITY = 1'b0;
    defparam \CPU/add_33/i29 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_33/i28  (.I0(n1533), .I1(\CPU/rs1[27] ), .CI(n668), 
            .O(n665), .CO(n666)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(131)
    defparam \CPU/add_33/i28 .I0_POLARITY = 1'b0;
    defparam \CPU/add_33/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_33/i27  (.I0(n1535), .I1(\CPU/rs1[26] ), .CI(n670), 
            .O(n667), .CO(n668)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(131)
    defparam \CPU/add_33/i27 .I0_POLARITY = 1'b0;
    defparam \CPU/add_33/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_33/i26  (.I0(n1537), .I1(\CPU/rs1[25] ), .CI(n672), 
            .O(n669), .CO(n670)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(131)
    defparam \CPU/add_33/i26 .I0_POLARITY = 1'b0;
    defparam \CPU/add_33/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_33/i25  (.I0(n1539), .I1(\CPU/rs1[24] ), .CI(n674), 
            .O(n671), .CO(n672)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(131)
    defparam \CPU/add_33/i25 .I0_POLARITY = 1'b0;
    defparam \CPU/add_33/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_33/i24  (.I0(n1541), .I1(\CPU/rs1[23] ), .CI(n676), 
            .O(n673), .CO(n674)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(131)
    defparam \CPU/add_33/i24 .I0_POLARITY = 1'b0;
    defparam \CPU/add_33/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_33/i23  (.I0(n1543), .I1(\CPU/rs1[22] ), .CI(n678), 
            .O(n675), .CO(n676)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(131)
    defparam \CPU/add_33/i23 .I0_POLARITY = 1'b0;
    defparam \CPU/add_33/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_33/i22  (.I0(n1545), .I1(\CPU/rs1[21] ), .CI(n680), 
            .O(n677), .CO(n678)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(131)
    defparam \CPU/add_33/i22 .I0_POLARITY = 1'b0;
    defparam \CPU/add_33/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_33/i21  (.I0(n1547), .I1(\CPU/rs1[20] ), .CI(n682), 
            .O(n679), .CO(n680)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(131)
    defparam \CPU/add_33/i21 .I0_POLARITY = 1'b0;
    defparam \CPU/add_33/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_33/i20  (.I0(n1549), .I1(\CPU/rs1[19] ), .CI(n684), 
            .O(n681), .CO(n682)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(131)
    defparam \CPU/add_33/i20 .I0_POLARITY = 1'b0;
    defparam \CPU/add_33/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_33/i19  (.I0(n1551), .I1(\CPU/rs1[18] ), .CI(n686), 
            .O(n683), .CO(n684)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(131)
    defparam \CPU/add_33/i19 .I0_POLARITY = 1'b0;
    defparam \CPU/add_33/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_33/i18  (.I0(n1553), .I1(\CPU/rs1[17] ), .CI(n688), 
            .O(n685), .CO(n686)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(131)
    defparam \CPU/add_33/i18 .I0_POLARITY = 1'b0;
    defparam \CPU/add_33/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_33/i17  (.I0(n1555), .I1(\CPU/rs1[16] ), .CI(n690), 
            .O(n687), .CO(n688)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(131)
    defparam \CPU/add_33/i17 .I0_POLARITY = 1'b0;
    defparam \CPU/add_33/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_33/i16  (.I0(n1557), .I1(\CPU/rs1[15] ), .CI(n692), 
            .O(n689), .CO(n690)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(131)
    defparam \CPU/add_33/i16 .I0_POLARITY = 1'b0;
    defparam \CPU/add_33/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_33/i15  (.I0(n1559), .I1(\CPU/rs1[14] ), .CI(n694), 
            .O(n691), .CO(n692)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(131)
    defparam \CPU/add_33/i15 .I0_POLARITY = 1'b0;
    defparam \CPU/add_33/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_33/i14  (.I0(n1561), .I1(\CPU/rs1[13] ), .CI(n696), 
            .O(n693), .CO(n694)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(131)
    defparam \CPU/add_33/i14 .I0_POLARITY = 1'b0;
    defparam \CPU/add_33/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_33/i13  (.I0(n1563), .I1(\CPU/rs1[12] ), .CI(n698), 
            .O(n695), .CO(n696)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(131)
    defparam \CPU/add_33/i13 .I0_POLARITY = 1'b0;
    defparam \CPU/add_33/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_33/i12  (.I0(n1565), .I1(\CPU/rs1[11] ), .CI(n700), 
            .O(n697), .CO(n698)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(131)
    defparam \CPU/add_33/i12 .I0_POLARITY = 1'b0;
    defparam \CPU/add_33/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_33/i11  (.I0(n1567), .I1(\CPU/rs1[10] ), .CI(n702), 
            .O(n699), .CO(n700)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(131)
    defparam \CPU/add_33/i11 .I0_POLARITY = 1'b0;
    defparam \CPU/add_33/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_33/i10  (.I0(n1569), .I1(\CPU/rs1[9] ), .CI(n704), 
            .O(n701), .CO(n702)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(131)
    defparam \CPU/add_33/i10 .I0_POLARITY = 1'b0;
    defparam \CPU/add_33/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_33/i9  (.I0(n1571), .I1(\CPU/rs1[8] ), .CI(n706), 
            .O(n703), .CO(n704)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(131)
    defparam \CPU/add_33/i9 .I0_POLARITY = 1'b0;
    defparam \CPU/add_33/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_33/i8  (.I0(n1573), .I1(\CPU/rs1[7] ), .CI(n708), 
            .O(n705), .CO(n706)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(131)
    defparam \CPU/add_33/i8 .I0_POLARITY = 1'b0;
    defparam \CPU/add_33/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_33/i7  (.I0(n1575), .I1(\CPU/rs1[6] ), .CI(n710), 
            .O(n707), .CO(n708)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(131)
    defparam \CPU/add_33/i7 .I0_POLARITY = 1'b0;
    defparam \CPU/add_33/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_33/i6  (.I0(n1577), .I1(\CPU/rs1[5] ), .CI(n712), 
            .O(n709), .CO(n710)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(131)
    defparam \CPU/add_33/i6 .I0_POLARITY = 1'b0;
    defparam \CPU/add_33/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_33/i5  (.I0(n1579), .I1(\CPU/rs1[4] ), .CI(n714), 
            .O(n711), .CO(n712)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(131)
    defparam \CPU/add_33/i5 .I0_POLARITY = 1'b0;
    defparam \CPU/add_33/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_33/i4  (.I0(n1581), .I1(\CPU/rs1[3] ), .CI(n716), 
            .O(n713), .CO(n714)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(131)
    defparam \CPU/add_33/i4 .I0_POLARITY = 1'b0;
    defparam \CPU/add_33/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_33/i3  (.I0(n1583), .I1(\CPU/rs1[2] ), .CI(n718), 
            .O(n715), .CO(n716)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(131)
    defparam \CPU/add_33/i3 .I0_POLARITY = 1'b0;
    defparam \CPU/add_33/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_33/i2  (.I0(n1585), .I1(\CPU/rs1[1] ), .CI(n7), .O(n717), 
            .CO(n718)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(131)
    defparam \CPU/add_33/i2 .I0_POLARITY = 1'b0;
    defparam \CPU/add_33/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_30/i32  (.I0(\CPU/rs1[31] ), .I1(n1525), .CI(n721), 
            .O(n719)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(127)
    defparam \CPU/add_30/i32 .I0_POLARITY = 1'b1;
    defparam \CPU/add_30/i32 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_30/i31  (.I0(\CPU/rs1[30] ), .I1(n1527), .CI(n723), 
            .O(n720), .CO(n721)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(127)
    defparam \CPU/add_30/i31 .I0_POLARITY = 1'b1;
    defparam \CPU/add_30/i31 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_30/i30  (.I0(\CPU/rs1[29] ), .I1(n1529), .CI(n725), 
            .O(n722), .CO(n723)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(127)
    defparam \CPU/add_30/i30 .I0_POLARITY = 1'b1;
    defparam \CPU/add_30/i30 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_30/i29  (.I0(\CPU/rs1[28] ), .I1(n1531), .CI(n727), 
            .O(n724), .CO(n725)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(127)
    defparam \CPU/add_30/i29 .I0_POLARITY = 1'b1;
    defparam \CPU/add_30/i29 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_30/i28  (.I0(\CPU/rs1[27] ), .I1(n1533), .CI(n729), 
            .O(n726), .CO(n727)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(127)
    defparam \CPU/add_30/i28 .I0_POLARITY = 1'b1;
    defparam \CPU/add_30/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_30/i27  (.I0(\CPU/rs1[26] ), .I1(n1535), .CI(n731), 
            .O(n728), .CO(n729)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(127)
    defparam \CPU/add_30/i27 .I0_POLARITY = 1'b1;
    defparam \CPU/add_30/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_30/i26  (.I0(\CPU/rs1[25] ), .I1(n1537), .CI(n733), 
            .O(n730), .CO(n731)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(127)
    defparam \CPU/add_30/i26 .I0_POLARITY = 1'b1;
    defparam \CPU/add_30/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_30/i25  (.I0(\CPU/rs1[24] ), .I1(n1539), .CI(n735), 
            .O(n732), .CO(n733)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(127)
    defparam \CPU/add_30/i25 .I0_POLARITY = 1'b1;
    defparam \CPU/add_30/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_30/i24  (.I0(\CPU/rs1[23] ), .I1(n1541), .CI(n737), 
            .O(n734), .CO(n735)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(127)
    defparam \CPU/add_30/i24 .I0_POLARITY = 1'b1;
    defparam \CPU/add_30/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_30/i23  (.I0(\CPU/rs1[22] ), .I1(n1543), .CI(n739), 
            .O(n736), .CO(n737)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(127)
    defparam \CPU/add_30/i23 .I0_POLARITY = 1'b1;
    defparam \CPU/add_30/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_30/i22  (.I0(\CPU/rs1[21] ), .I1(n1545), .CI(n741), 
            .O(n738), .CO(n739)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(127)
    defparam \CPU/add_30/i22 .I0_POLARITY = 1'b1;
    defparam \CPU/add_30/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_30/i21  (.I0(\CPU/rs1[20] ), .I1(n1547), .CI(n743), 
            .O(n740), .CO(n741)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(127)
    defparam \CPU/add_30/i21 .I0_POLARITY = 1'b1;
    defparam \CPU/add_30/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_30/i20  (.I0(\CPU/rs1[19] ), .I1(n1549), .CI(n745), 
            .O(n742), .CO(n743)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(127)
    defparam \CPU/add_30/i20 .I0_POLARITY = 1'b1;
    defparam \CPU/add_30/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_30/i19  (.I0(\CPU/rs1[18] ), .I1(n1551), .CI(n747), 
            .O(n744), .CO(n745)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(127)
    defparam \CPU/add_30/i19 .I0_POLARITY = 1'b1;
    defparam \CPU/add_30/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_30/i18  (.I0(\CPU/rs1[17] ), .I1(n1553), .CI(n749), 
            .O(n746), .CO(n747)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(127)
    defparam \CPU/add_30/i18 .I0_POLARITY = 1'b1;
    defparam \CPU/add_30/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_30/i17  (.I0(\CPU/rs1[16] ), .I1(n1555), .CI(n751), 
            .O(n748), .CO(n749)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(127)
    defparam \CPU/add_30/i17 .I0_POLARITY = 1'b1;
    defparam \CPU/add_30/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_30/i16  (.I0(\CPU/rs1[15] ), .I1(n1557), .CI(n753), 
            .O(n750), .CO(n751)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(127)
    defparam \CPU/add_30/i16 .I0_POLARITY = 1'b1;
    defparam \CPU/add_30/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_30/i15  (.I0(\CPU/rs1[14] ), .I1(n1559), .CI(n755), 
            .O(n752), .CO(n753)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(127)
    defparam \CPU/add_30/i15 .I0_POLARITY = 1'b1;
    defparam \CPU/add_30/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_30/i14  (.I0(\CPU/rs1[13] ), .I1(n1561), .CI(n757), 
            .O(n754), .CO(n755)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(127)
    defparam \CPU/add_30/i14 .I0_POLARITY = 1'b1;
    defparam \CPU/add_30/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_30/i13  (.I0(\CPU/rs1[12] ), .I1(n1563), .CI(n759), 
            .O(n756), .CO(n757)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(127)
    defparam \CPU/add_30/i13 .I0_POLARITY = 1'b1;
    defparam \CPU/add_30/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_30/i12  (.I0(\CPU/rs1[11] ), .I1(n1565), .CI(n761), 
            .O(n758), .CO(n759)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(127)
    defparam \CPU/add_30/i12 .I0_POLARITY = 1'b1;
    defparam \CPU/add_30/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_30/i11  (.I0(\CPU/rs1[10] ), .I1(n1567), .CI(n763), 
            .O(n760), .CO(n761)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(127)
    defparam \CPU/add_30/i11 .I0_POLARITY = 1'b1;
    defparam \CPU/add_30/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_30/i10  (.I0(\CPU/rs1[9] ), .I1(n1569), .CI(n765), 
            .O(n762), .CO(n763)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(127)
    defparam \CPU/add_30/i10 .I0_POLARITY = 1'b1;
    defparam \CPU/add_30/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_30/i9  (.I0(\CPU/rs1[8] ), .I1(n1571), .CI(n767), 
            .O(n764), .CO(n765)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(127)
    defparam \CPU/add_30/i9 .I0_POLARITY = 1'b1;
    defparam \CPU/add_30/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_30/i8  (.I0(\CPU/rs1[7] ), .I1(n1573), .CI(n769), 
            .O(n766), .CO(n767)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(127)
    defparam \CPU/add_30/i8 .I0_POLARITY = 1'b1;
    defparam \CPU/add_30/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_30/i7  (.I0(\CPU/rs1[6] ), .I1(n1575), .CI(n771), 
            .O(n768), .CO(n769)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(127)
    defparam \CPU/add_30/i7 .I0_POLARITY = 1'b1;
    defparam \CPU/add_30/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_30/i6  (.I0(\CPU/rs1[5] ), .I1(n1577), .CI(n773), 
            .O(n770), .CO(n771)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(127)
    defparam \CPU/add_30/i6 .I0_POLARITY = 1'b1;
    defparam \CPU/add_30/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_30/i5  (.I0(\CPU/rs1[4] ), .I1(n1579), .CI(n775), 
            .O(n772), .CO(n773)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(127)
    defparam \CPU/add_30/i5 .I0_POLARITY = 1'b1;
    defparam \CPU/add_30/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_30/i4  (.I0(\CPU/rs1[3] ), .I1(n1581), .CI(n777), 
            .O(n774), .CO(n775)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(127)
    defparam \CPU/add_30/i4 .I0_POLARITY = 1'b1;
    defparam \CPU/add_30/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_30/i3  (.I0(\CPU/rs1[2] ), .I1(n1583), .CI(n779), 
            .O(n776), .CO(n777)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(127)
    defparam \CPU/add_30/i3 .I0_POLARITY = 1'b1;
    defparam \CPU/add_30/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_30/i2  (.I0(\CPU/rs1[1] ), .I1(n1585), .CI(n781), 
            .O(n778), .CO(n779)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(127)
    defparam \CPU/add_30/i2 .I0_POLARITY = 1'b1;
    defparam \CPU/add_30/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \CPU/add_30/i1  (.I0(\CPU/rs1[0] ), .I1(n1587), .CI(1'b0), 
            .O(n780), .CO(n781)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(127)
    defparam \CPU/add_30/i1 .I0_POLARITY = 1'b1;
    defparam \CPU/add_30/i1 .I1_POLARITY = 1'b1;
    EFX_RAM_5K \RAM/MEM__D$c12  (.WCLK(\clk~O ), .RCLK(\clk~O ), .WCLKE(1'b1), 
            .WE(\RAM/n116 ), .RE(n107), .WDATA({\mem_wdata[24] }), .WADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RDATA({\RAM_rdata[24] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h1102050461089300020000A4A008204001404004042926800002890006800008, INIT_1=256'h0000000000006D10EA12820810102638C00A00C0280291930250142299268020, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/bram/bram.v(12)
    defparam \RAM/MEM__D$c12 .READ_WIDTH = 1;
    defparam \RAM/MEM__D$c12 .WRITE_WIDTH = 1;
    defparam \RAM/MEM__D$c12 .WCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$c12 .WCLKE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$c12 .WE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$c12 .RCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$c12 .RE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$c12 .INIT_0 = 256'h1102050461089300020000A4A008204001404004042926800002890006800008;
    defparam \RAM/MEM__D$c12 .INIT_1 = 256'h0000000000006D10EA12820810102638C00A00C0280291930250142299268020;
    defparam \RAM/MEM__D$c12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$c12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$c12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$c12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$c12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$c12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$c12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$c12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$c12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$c12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$c12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$c12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$c12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$c12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$c12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$c12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$c12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$c12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$c12 .OUTPUT_REG = 1'b0;
    defparam \RAM/MEM__D$c12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \CPU/registerFile__D$1  (.WCLK(\clk~O ), .RCLK(\clk~O ), 
            .WCLKE(\CPU/writeBack ), .WE(\CPU/not_equal_22/n9 ), .RE(\CPU/n3447 ), 
            .WDATA({\CPU/writeBackData[31] , \CPU/writeBackData[30] , \CPU/writeBackData[29] , 
            \CPU/writeBackData[28] , \CPU/writeBackData[27] , \CPU/writeBackData[26] , 
            \CPU/writeBackData[25] , \CPU/writeBackData[24] , \CPU/writeBackData[23] , 
            \CPU/writeBackData[22] , \CPU/writeBackData[21] , \CPU/writeBackData[20] , 
            \CPU/writeBackData[19] , \CPU/writeBackData[18] , \CPU/writeBackData[17] , 
            \CPU/writeBackData[16] }), .WADDR({3'b000, \CPU/instr[11] , 
            \CPU/instr[10] , \CPU/instr[9] , \CPU/instr[8] , \CPU/instr[7] }), 
            .RADDR({3'b000, \mem_rdata[19] , \mem_rdata[18] , \mem_rdata[17] , 
            \mem_rdata[16] , \mem_rdata[15] }), .RDATA({\CPU/rs1[31] , 
            \CPU/rs1[30] , \CPU/rs1[29] , \CPU/rs1[28] , \CPU/rs1[27] , 
            \CPU/rs1[26] , \CPU/rs1[25] , \CPU/rs1[24] , \CPU/rs1[23] , 
            \CPU/rs1[22] , \CPU/rs1[21] , \CPU/rs1[20] , \CPU/rs1[19] , 
            \CPU/rs1[18] , \CPU/rs1[17] , \CPU/rs1[16] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=16, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(100)
    defparam \CPU/registerFile__D$1 .READ_WIDTH = 16;
    defparam \CPU/registerFile__D$1 .WRITE_WIDTH = 16;
    defparam \CPU/registerFile__D$1 .WCLK_POLARITY = 1'b1;
    defparam \CPU/registerFile__D$1 .WCLKE_POLARITY = 1'b1;
    defparam \CPU/registerFile__D$1 .WE_POLARITY = 1'b1;
    defparam \CPU/registerFile__D$1 .RCLK_POLARITY = 1'b1;
    defparam \CPU/registerFile__D$1 .RE_POLARITY = 1'b1;
    defparam \CPU/registerFile__D$1 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$1 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$1 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$1 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$1 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$1 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$1 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$1 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$1 .OUTPUT_REG = 1'b0;
    defparam \CPU/registerFile__D$1 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \CPU/registerFile__D$2  (.WCLK(\clk~O ), .RCLK(\clk~O ), 
            .WCLKE(\CPU/writeBack ), .WE(\CPU/not_equal_22/n9 ), .RE(\CPU/n3447 ), 
            .WDATA({\CPU/writeBackData[15] , \CPU/writeBackData[14] , \CPU/writeBackData[13] , 
            \CPU/writeBackData[12] , \CPU/writeBackData[11] , \CPU/writeBackData[10] , 
            \CPU/writeBackData[9] , \CPU/writeBackData[8] , \CPU/writeBackData[7] , 
            \CPU/writeBackData[6] , \CPU/writeBackData[5] , \CPU/writeBackData[4] , 
            \CPU/writeBackData[3] , \CPU/writeBackData[2] , \CPU/writeBackData[1] , 
            \CPU/writeBackData[0] }), .WADDR({3'b000, \CPU/instr[11] , 
            \CPU/instr[10] , \CPU/instr[9] , \CPU/instr[8] , \CPU/instr[7] }), 
            .RADDR({3'b000, \mem_rdata[19] , \mem_rdata[18] , \mem_rdata[17] , 
            \mem_rdata[16] , \mem_rdata[15] }), .RDATA({\CPU/rs1[15] , 
            \CPU/rs1[14] , \CPU/rs1[13] , \CPU/rs1[12] , \CPU/rs1[11] , 
            \CPU/rs1[10] , \CPU/rs1[9] , \CPU/rs1[8] , \CPU/rs1[7] , 
            \CPU/rs1[6] , \CPU/rs1[5] , \CPU/rs1[4] , \CPU/rs1[3] , 
            \CPU/rs1[2] , \CPU/rs1[1] , \CPU/rs1[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=16, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(100)
    defparam \CPU/registerFile__D$2 .READ_WIDTH = 16;
    defparam \CPU/registerFile__D$2 .WRITE_WIDTH = 16;
    defparam \CPU/registerFile__D$2 .WCLK_POLARITY = 1'b1;
    defparam \CPU/registerFile__D$2 .WCLKE_POLARITY = 1'b1;
    defparam \CPU/registerFile__D$2 .WE_POLARITY = 1'b1;
    defparam \CPU/registerFile__D$2 .RCLK_POLARITY = 1'b1;
    defparam \CPU/registerFile__D$2 .RE_POLARITY = 1'b1;
    defparam \CPU/registerFile__D$2 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$2 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$2 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$2 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$2 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$2 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$2 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$2 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$2 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$2 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$2 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$2 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$2 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$2 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$2 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$2 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$2 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$2 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$2 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$2 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile__D$2 .OUTPUT_REG = 1'b0;
    defparam \CPU/registerFile__D$2 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \CPU/registerFile_2__D$2  (.WCLK(\clk~O ), .RCLK(\clk~O ), 
            .WCLKE(\CPU/writeBack ), .WE(\CPU/not_equal_22/n9 ), .RE(\CPU/n3447 ), 
            .WDATA({\CPU/writeBackData[15] , \CPU/writeBackData[14] , \CPU/writeBackData[13] , 
            \CPU/writeBackData[12] , \CPU/writeBackData[11] , \CPU/writeBackData[10] , 
            \CPU/writeBackData[9] , \CPU/writeBackData[8] , \CPU/writeBackData[7] , 
            \CPU/writeBackData[6] , \CPU/writeBackData[5] , \CPU/writeBackData[4] , 
            \CPU/writeBackData[3] , \CPU/writeBackData[2] , \CPU/writeBackData[1] , 
            \CPU/writeBackData[0] }), .WADDR({3'b000, \CPU/instr[11] , 
            \CPU/instr[10] , \CPU/instr[9] , \CPU/instr[8] , \CPU/instr[7] }), 
            .RADDR({3'b000, \mem_rdata[24] , \mem_rdata[23] , \mem_rdata[22] , 
            \mem_rdata[21] , \mem_rdata[20] }), .RDATA({\CPU/rs2[15] , 
            \CPU/rs2[14] , \CPU/rs2[13] , \CPU/rs2[12] , \CPU/rs2[11] , 
            \CPU/rs2[10] , \CPU/rs2[9] , \CPU/rs2[8] , \mem_wdata[7] , 
            \mem_wdata[6] , \mem_wdata[5] , \mem_wdata[4] , \mem_wdata[3] , 
            \mem_wdata[2] , \mem_wdata[1] , \mem_wdata[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=16, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(100)
    defparam \CPU/registerFile_2__D$2 .READ_WIDTH = 16;
    defparam \CPU/registerFile_2__D$2 .WRITE_WIDTH = 16;
    defparam \CPU/registerFile_2__D$2 .WCLK_POLARITY = 1'b1;
    defparam \CPU/registerFile_2__D$2 .WCLKE_POLARITY = 1'b1;
    defparam \CPU/registerFile_2__D$2 .WE_POLARITY = 1'b1;
    defparam \CPU/registerFile_2__D$2 .RCLK_POLARITY = 1'b1;
    defparam \CPU/registerFile_2__D$2 .RE_POLARITY = 1'b1;
    defparam \CPU/registerFile_2__D$2 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$2 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$2 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$2 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$2 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$2 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$2 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$2 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$2 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$2 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$2 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$2 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$2 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$2 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$2 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$2 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$2 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$2 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$2 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$2 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$2 .OUTPUT_REG = 1'b0;
    defparam \CPU/registerFile_2__D$2 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \CPU/registerFile_2__D$1  (.WCLK(\clk~O ), .RCLK(\clk~O ), 
            .WCLKE(\CPU/writeBack ), .WE(\CPU/not_equal_22/n9 ), .RE(\CPU/n3447 ), 
            .WDATA({\CPU/writeBackData[31] , \CPU/writeBackData[30] , \CPU/writeBackData[29] , 
            \CPU/writeBackData[28] , \CPU/writeBackData[27] , \CPU/writeBackData[26] , 
            \CPU/writeBackData[25] , \CPU/writeBackData[24] , \CPU/writeBackData[23] , 
            \CPU/writeBackData[22] , \CPU/writeBackData[21] , \CPU/writeBackData[20] , 
            \CPU/writeBackData[19] , \CPU/writeBackData[18] , \CPU/writeBackData[17] , 
            \CPU/writeBackData[16] }), .WADDR({3'b000, \CPU/instr[11] , 
            \CPU/instr[10] , \CPU/instr[9] , \CPU/instr[8] , \CPU/instr[7] }), 
            .RADDR({3'b000, \mem_rdata[24] , \mem_rdata[23] , \mem_rdata[22] , 
            \mem_rdata[21] , \mem_rdata[20] }), .RDATA({\CPU/rs2[31] , 
            \CPU/rs2[30] , \CPU/rs2[29] , \CPU/rs2[28] , \CPU/rs2[27] , 
            \CPU/rs2[26] , \CPU/rs2[25] , \CPU/rs2[24] , \CPU/rs2[23] , 
            \CPU/rs2[22] , \CPU/rs2[21] , \CPU/rs2[20] , \CPU/rs2[19] , 
            \CPU/rs2[18] , \CPU/rs2[17] , \CPU/rs2[16] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=16, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(100)
    defparam \CPU/registerFile_2__D$1 .READ_WIDTH = 16;
    defparam \CPU/registerFile_2__D$1 .WRITE_WIDTH = 16;
    defparam \CPU/registerFile_2__D$1 .WCLK_POLARITY = 1'b1;
    defparam \CPU/registerFile_2__D$1 .WCLKE_POLARITY = 1'b1;
    defparam \CPU/registerFile_2__D$1 .WE_POLARITY = 1'b1;
    defparam \CPU/registerFile_2__D$1 .RCLK_POLARITY = 1'b1;
    defparam \CPU/registerFile_2__D$1 .RE_POLARITY = 1'b1;
    defparam \CPU/registerFile_2__D$1 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$1 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$1 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$1 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$1 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$1 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$1 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$1 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CPU/registerFile_2__D$1 .OUTPUT_REG = 1'b0;
    defparam \CPU/registerFile_2__D$1 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \RAM/MEM__D$2b12  (.WCLK(\clk~O ), .RCLK(\clk~O ), .WCLKE(1'b1), 
            .WE(\RAM/n104 ), .RE(n107), .WDATA({\mem_wdata[2] }), .WADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RDATA({\RAM_rdata[2] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'hC040600638C0083604006202129514A223229228060C10C0001C70E81B70403F, INIT_1=256'h0000000000004201E83CDE408020031C7007007007000080002006108010C040, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/bram/bram.v(12)
    defparam \RAM/MEM__D$2b12 .READ_WIDTH = 1;
    defparam \RAM/MEM__D$2b12 .WRITE_WIDTH = 1;
    defparam \RAM/MEM__D$2b12 .WCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$2b12 .WCLKE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$2b12 .WE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$2b12 .RCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$2b12 .RE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$2b12 .INIT_0 = 256'hC040600638C0083604006202129514A223229228060C10C0001C70E81B70403F;
    defparam \RAM/MEM__D$2b12 .INIT_1 = 256'h0000000000004201E83CDE408020031C7007007007000080002006108010C040;
    defparam \RAM/MEM__D$2b12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2b12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2b12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2b12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2b12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2b12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2b12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2b12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2b12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2b12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2b12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2b12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2b12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2b12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2b12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2b12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2b12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2b12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2b12 .OUTPUT_REG = 1'b0;
    defparam \RAM/MEM__D$2b12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \RAM/MEM__D$b1b2  (.WCLK(\clk~O ), .RCLK(\clk~O ), .WCLKE(1'b1), 
            .WE(\RAM/n112 ), .RE(n107), .WDATA({\mem_wdata[16] }), .WADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RDATA({\RAM_rdata[16] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h392492590410F7807B99183DE96AAB5454956DC72851EE3FF9F18514408903E0, INIT_1=256'h0000000000018614EA97DDAB755EC8C30D50D50D50D52A2003DC91EC31EE07BC, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/bram/bram.v(12)
    defparam \RAM/MEM__D$b1b2 .READ_WIDTH = 1;
    defparam \RAM/MEM__D$b1b2 .WRITE_WIDTH = 1;
    defparam \RAM/MEM__D$b1b2 .WCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b1b2 .WCLKE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b1b2 .WE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b1b2 .RCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b1b2 .RE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b1b2 .INIT_0 = 256'h392492590410F7807B99183DE96AAB5454956DC72851EE3FF9F18514408903E0;
    defparam \RAM/MEM__D$b1b2 .INIT_1 = 256'h0000000000018614EA97DDAB755EC8C30D50D50D50D52A2003DC91EC31EE07BC;
    defparam \RAM/MEM__D$b1b2 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b1b2 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b1b2 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b1b2 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b1b2 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b1b2 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b1b2 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b1b2 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b1b2 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b1b2 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b1b2 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b1b2 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b1b2 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b1b2 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b1b2 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b1b2 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b1b2 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b1b2 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b1b2 .OUTPUT_REG = 1'b0;
    defparam \RAM/MEM__D$b1b2 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \RAM/MEM__D$d12  (.WCLK(\clk~O ), .RCLK(\clk~O ), .WCLKE(1'b1), 
            .WE(\RAM/n116 ), .RE(n107), .WDATA({\mem_wdata[25] }), .WADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RDATA({\RAM_rdata[25] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h97FC41A40036E401CB86C73904004019004841473481C80007222815B606AE40, INIT_1=256'h000000000001E425B43434AC400C820062E62E02E22E0C6403DC7C21D1C82CBB, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/bram/bram.v(12)
    defparam \RAM/MEM__D$d12 .READ_WIDTH = 1;
    defparam \RAM/MEM__D$d12 .WRITE_WIDTH = 1;
    defparam \RAM/MEM__D$d12 .WCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$d12 .WCLKE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$d12 .WE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$d12 .RCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$d12 .RE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$d12 .INIT_0 = 256'h97FC41A40036E401CB86C73904004019004841473481C80007222815B606AE40;
    defparam \RAM/MEM__D$d12 .INIT_1 = 256'h000000000001E425B43434AC400C820062E62E02E22E0C6403DC7C21D1C82CBB;
    defparam \RAM/MEM__D$d12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$d12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$d12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$d12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$d12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$d12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$d12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$d12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$d12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$d12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$d12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$d12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$d12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$d12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$d12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$d12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$d12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$d12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$d12 .OUTPUT_REG = 1'b0;
    defparam \RAM/MEM__D$d12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \RAM/MEM__D$12b12  (.WCLK(\clk~O ), .RCLK(\clk~O ), .WCLKE(1'b1), 
            .WE(\RAM/n108 ), .RE(n107), .WDATA({\mem_wdata[10] }), .WADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RDATA({\RAM_rdata[10] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h3F9B9DF9C72FE2C9F11F9DF8FEFDF7EFFEEFF78218F3C43FFFC2CB9BE4CFBF80, INIT_1=256'h0000000000015B9B0BE3CEAD404B7CE38FB8FB8FB8FBFF7F378879FF7FC43F13, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/bram/bram.v(12)
    defparam \RAM/MEM__D$12b12 .READ_WIDTH = 1;
    defparam \RAM/MEM__D$12b12 .WRITE_WIDTH = 1;
    defparam \RAM/MEM__D$12b12 .WCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$12b12 .WCLKE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$12b12 .WE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$12b12 .RCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$12b12 .RE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$12b12 .INIT_0 = 256'h3F9B9DF9C72FE2C9F11F9DF8FEFDF7EFFEEFF78218F3C43FFFC2CB9BE4CFBF80;
    defparam \RAM/MEM__D$12b12 .INIT_1 = 256'h0000000000015B9B0BE3CEAD404B7CE38FB8FB8FB8FBFF7F378879FF7FC43F13;
    defparam \RAM/MEM__D$12b12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12b12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12b12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12b12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12b12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12b12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12b12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12b12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12b12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12b12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12b12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12b12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12b12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12b12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12b12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12b12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12b12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12b12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12b12 .OUTPUT_REG = 1'b0;
    defparam \RAM/MEM__D$12b12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \RAM/MEM__D$b2  (.WCLK(\clk~O ), .RCLK(\clk~O ), .WCLKE(1'b1), 
            .WE(\RAM/n104 ), .RE(n107), .WDATA({\mem_wdata[0] }), .WADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RDATA({\RAM_rdata[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_1=256'h000000000001041ECBCF0DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/bram/bram.v(12)
    defparam \RAM/MEM__D$b2 .READ_WIDTH = 1;
    defparam \RAM/MEM__D$b2 .WRITE_WIDTH = 1;
    defparam \RAM/MEM__D$b2 .WCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b2 .WCLKE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b2 .WE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b2 .RCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b2 .RE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b2 .INIT_0 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \RAM/MEM__D$b2 .INIT_1 = 256'h000000000001041ECBCF0DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \RAM/MEM__D$b2 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b2 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b2 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b2 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b2 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b2 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b2 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b2 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b2 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b2 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b2 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b2 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b2 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b2 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b2 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b2 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b2 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b2 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b2 .OUTPUT_REG = 1'b0;
    defparam \RAM/MEM__D$b2 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \RAM/MEM__D$1b2  (.WCLK(\clk~O ), .RCLK(\clk~O ), .WCLKE(1'b1), 
            .WE(\RAM/n108 ), .RE(n107), .WDATA({\mem_wdata[8] }), .WADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RDATA({\RAM_rdata[8] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h3D9A9D69C72A14C90A0D9C8576FDF7EEBE6EF6441870283FFC22CB9BE4CFBC53, INIT_1=256'h000000000000F19F0BE2050930136CE38DB8DB8DB8DBB734005059FF382830A3, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/bram/bram.v(12)
    defparam \RAM/MEM__D$1b2 .READ_WIDTH = 1;
    defparam \RAM/MEM__D$1b2 .WRITE_WIDTH = 1;
    defparam \RAM/MEM__D$1b2 .WCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$1b2 .WCLKE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$1b2 .WE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$1b2 .RCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$1b2 .RE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$1b2 .INIT_0 = 256'h3D9A9D69C72A14C90A0D9C8576FDF7EEBE6EF6441870283FFC22CB9BE4CFBC53;
    defparam \RAM/MEM__D$1b2 .INIT_1 = 256'h000000000000F19F0BE2050930136CE38DB8DB8DB8DBB734005059FF382830A3;
    defparam \RAM/MEM__D$1b2 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$1b2 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$1b2 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$1b2 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$1b2 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$1b2 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$1b2 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$1b2 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$1b2 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$1b2 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$1b2 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$1b2 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$1b2 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$1b2 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$1b2 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$1b2 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$1b2 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$1b2 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$1b2 .OUTPUT_REG = 1'b0;
    defparam \RAM/MEM__D$1b2 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \RAM/MEM__D$e12  (.WCLK(\clk~O ), .RCLK(\clk~O ), .WCLKE(1'b1), 
            .WE(\RAM/n116 ), .RE(n107), .WDATA({\mem_wdata[26] }), .WADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RDATA({\RAM_rdata[26] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h879B45A4511F1021881685C42D2A694D44C54C4030AA200006320841B226EC40, INIT_1=256'h0000000000014514AA12F32C4010B428A2AE2A82AC2AD9780400F8035E202887, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/bram/bram.v(12)
    defparam \RAM/MEM__D$e12 .READ_WIDTH = 1;
    defparam \RAM/MEM__D$e12 .WRITE_WIDTH = 1;
    defparam \RAM/MEM__D$e12 .WCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$e12 .WCLKE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$e12 .WE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$e12 .RCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$e12 .RE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$e12 .INIT_0 = 256'h879B45A4511F1021881685C42D2A694D44C54C4030AA200006320841B226EC40;
    defparam \RAM/MEM__D$e12 .INIT_1 = 256'h0000000000014514AA12F32C4010B428A2AE2A82AC2AD9780400F8035E202887;
    defparam \RAM/MEM__D$e12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$e12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$e12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$e12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$e12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$e12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$e12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$e12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$e12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$e12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$e12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$e12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$e12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$e12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$e12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$e12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$e12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$e12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$e12 .OUTPUT_REG = 1'b0;
    defparam \RAM/MEM__D$e12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \RAM/MEM__D$b12b12  (.WCLK(\clk~O ), .RCLK(\clk~O ), .WCLKE(1'b1), 
            .WE(\RAM/n112 ), .RE(n107), .WDATA({\mem_wdata[18] }), .WADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RDATA({\RAM_rdata[18] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h3FBF97F9451F0081801F9DC06D6AEB5D54956C0038F2003FFE118515E08FAC00, INIT_1=256'h0000000000014E04848725AA0002FCE38FD8FD8FD8FDFB7FFC00F9EF7E002807, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/bram/bram.v(12)
    defparam \RAM/MEM__D$b12b12 .READ_WIDTH = 1;
    defparam \RAM/MEM__D$b12b12 .WRITE_WIDTH = 1;
    defparam \RAM/MEM__D$b12b12 .WCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b12b12 .WCLKE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b12b12 .WE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b12b12 .RCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b12b12 .RE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b12b12 .INIT_0 = 256'h3FBF97F9451F0081801F9DC06D6AEB5D54956C0038F2003FFE118515E08FAC00;
    defparam \RAM/MEM__D$b12b12 .INIT_1 = 256'h0000000000014E04848725AA0002FCE38FD8FD8FD8FDFB7FFC00F9EF7E002807;
    defparam \RAM/MEM__D$b12b12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12b12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12b12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12b12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12b12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12b12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12b12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12b12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12b12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12b12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12b12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12b12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12b12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12b12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12b12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12b12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12b12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12b12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12b12 .OUTPUT_REG = 1'b0;
    defparam \RAM/MEM__D$b12b12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \RAM/MEM__D$f12  (.WCLK(\clk~O ), .RCLK(\clk~O ), .WCLKE(1'b1), 
            .WE(\RAM/n116 ), .RE(n107), .WDATA({\mem_wdata[27] }), .WADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RDATA({\RAM_rdata[27] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h07BF45A0710F10058816C5C4040040090040004030A2200006320805A026AC60, INIT_1=256'h00000000000004044012482C4000B420828828E28C28D9780440FC035E202887, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/bram/bram.v(12)
    defparam \RAM/MEM__D$f12 .READ_WIDTH = 1;
    defparam \RAM/MEM__D$f12 .WRITE_WIDTH = 1;
    defparam \RAM/MEM__D$f12 .WCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$f12 .WCLKE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$f12 .WE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$f12 .RCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$f12 .RE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$f12 .INIT_0 = 256'h07BF45A0710F10058816C5C4040040090040004030A2200006320805A026AC60;
    defparam \RAM/MEM__D$f12 .INIT_1 = 256'h00000000000004044012482C4000B420828828E28C28D9780440FC035E202887;
    defparam \RAM/MEM__D$f12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$f12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$f12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$f12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$f12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$f12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$f12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$f12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$f12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$f12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$f12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$f12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$f12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$f12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$f12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$f12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$f12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$f12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$f12 .OUTPUT_REG = 1'b0;
    defparam \RAM/MEM__D$f12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \RAM/MEM__D$g12  (.WCLK(\clk~O ), .RCLK(\clk~O ), .WCLKE(1'b1), 
            .WE(\RAM/n116 ), .RE(n107), .WDATA({\mem_wdata[28] }), .WADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RDATA({\RAM_rdata[28] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h07B400A41084E0258816C5C42D2A694D44C5044030A2200006320815A0A6AC60, INIT_1=256'h00000000000060048010182640003420828A28828A28D1F80440FC235E2028BE, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/bram/bram.v(12)
    defparam \RAM/MEM__D$g12 .READ_WIDTH = 1;
    defparam \RAM/MEM__D$g12 .WRITE_WIDTH = 1;
    defparam \RAM/MEM__D$g12 .WCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$g12 .WCLKE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$g12 .WE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$g12 .RCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$g12 .RE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$g12 .INIT_0 = 256'h07B400A41084E0258816C5C42D2A694D44C5044030A2200006320815A0A6AC60;
    defparam \RAM/MEM__D$g12 .INIT_1 = 256'h00000000000060048010182640003420828A28828A28D1F80440FC235E2028BE;
    defparam \RAM/MEM__D$g12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$g12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$g12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$g12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$g12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$g12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$g12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$g12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$g12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$g12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$g12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$g12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$g12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$g12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$g12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$g12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$g12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$g12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$g12 .OUTPUT_REG = 1'b0;
    defparam \RAM/MEM__D$g12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \RAM/MEM__D$h12  (.WCLK(\clk~O ), .RCLK(\clk~O ), .WCLKE(1'b1), 
            .WE(\RAM/n116 ), .RE(n107), .WDATA({\mem_wdata[29] }), .WADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RDATA({\RAM_rdata[29] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h87BF44A4518F10258816C5C42D2A694D44C5044030A2200006300015A0A6AC40, INIT_1=256'h0000000000006F04801048244800B420828828A28828D1780440F8235E202887, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/bram/bram.v(12)
    defparam \RAM/MEM__D$h12 .READ_WIDTH = 1;
    defparam \RAM/MEM__D$h12 .WRITE_WIDTH = 1;
    defparam \RAM/MEM__D$h12 .WCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$h12 .WCLKE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$h12 .WE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$h12 .RCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$h12 .RE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$h12 .INIT_0 = 256'h87BF44A4518F10258816C5C42D2A694D44C5044030A2200006300015A0A6AC40;
    defparam \RAM/MEM__D$h12 .INIT_1 = 256'h0000000000006F04801048244800B420828828A28828D1780440F8235E202887;
    defparam \RAM/MEM__D$h12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$h12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$h12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$h12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$h12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$h12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$h12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$h12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$h12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$h12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$h12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$h12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$h12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$h12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$h12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$h12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$h12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$h12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$h12 .OUTPUT_REG = 1'b0;
    defparam \RAM/MEM__D$h12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \RAM/MEM__D$i12  (.WCLK(\clk~O ), .RCLK(\clk~O ), .WCLKE(1'b1), 
            .WE(\RAM/n116 ), .RE(n107), .WDATA({\mem_wdata[30] }), .WADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RDATA({\RAM_rdata[30] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h07BF04A0530F1005881685C42D6A694DC4C5044030A2200226300055A286AC40, INIT_1=256'h000000000001850E6140DC244000B420828A28A28A28D1780440F8235E202887, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/bram/bram.v(12)
    defparam \RAM/MEM__D$i12 .READ_WIDTH = 1;
    defparam \RAM/MEM__D$i12 .WRITE_WIDTH = 1;
    defparam \RAM/MEM__D$i12 .WCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$i12 .WCLKE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$i12 .WE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$i12 .RCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$i12 .RE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$i12 .INIT_0 = 256'h07BF04A0530F1005881685C42D6A694DC4C5044030A2200226300055A286AC40;
    defparam \RAM/MEM__D$i12 .INIT_1 = 256'h000000000001850E6140DC244000B420828A28A28A28D1780440F8235E202887;
    defparam \RAM/MEM__D$i12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$i12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$i12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$i12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$i12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$i12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$i12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$i12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$i12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$i12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$i12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$i12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$i12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$i12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$i12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$i12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$i12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$i12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$i12 .OUTPUT_REG = 1'b0;
    defparam \RAM/MEM__D$i12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \RAM/MEM__D$j1  (.WCLK(\clk~O ), .RCLK(\clk~O ), .WCLKE(1'b1), 
            .WE(\RAM/n116 ), .RE(n107), .WDATA({\mem_wdata[31] }), .WADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RDATA({\RAM_rdata[31] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h07BF04A0510F1005881685C4040040098040004030A2200006300005A006AC40, INIT_1=256'h0000000000000025342E06244000B420828A28A28A28D1780440F8035E202887, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/bram/bram.v(12)
    defparam \RAM/MEM__D$j1 .READ_WIDTH = 1;
    defparam \RAM/MEM__D$j1 .WRITE_WIDTH = 1;
    defparam \RAM/MEM__D$j1 .WCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$j1 .WCLKE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$j1 .WE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$j1 .RCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$j1 .RE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$j1 .INIT_0 = 256'h07BF04A0510F1005881685C4040040098040004030A2200006300005A006AC40;
    defparam \RAM/MEM__D$j1 .INIT_1 = 256'h0000000000000025342E06244000B420828A28A28A28D1780440F8035E202887;
    defparam \RAM/MEM__D$j1 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$j1 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$j1 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$j1 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$j1 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$j1 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$j1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$j1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$j1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$j1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$j1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$j1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$j1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$j1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$j1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$j1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$j1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$j1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$j1 .OUTPUT_REG = 1'b0;
    defparam \RAM/MEM__D$j1 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \RAM/MEM__D$b1212  (.WCLK(\clk~O ), .RCLK(\clk~O ), .WCLKE(1'b1), 
            .WE(\RAM/n112 ), .RE(n107), .WDATA({\mem_wdata[17] }), .WADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RDATA({\RAM_rdata[17] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h392413510410008000191800696AAB5454956C002040003FF811851440890020, INIT_1=256'h00000000000066317E287A046002C8C30D50D50D50D52A20000091EC30000004, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/bram/bram.v(12)
    defparam \RAM/MEM__D$b1212 .READ_WIDTH = 1;
    defparam \RAM/MEM__D$b1212 .WRITE_WIDTH = 1;
    defparam \RAM/MEM__D$b1212 .WCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b1212 .WCLKE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b1212 .WE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b1212 .RCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b1212 .RE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b1212 .INIT_0 = 256'h392413510410008000191800696AAB5454956C002040003FF811851440890020;
    defparam \RAM/MEM__D$b1212 .INIT_1 = 256'h00000000000066317E287A046002C8C30D50D50D50D52A20000091EC30000004;
    defparam \RAM/MEM__D$b1212 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b1212 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b1212 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b1212 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b1212 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b1212 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b1212 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b1212 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b1212 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b1212 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b1212 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b1212 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b1212 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b1212 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b1212 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b1212 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b1212 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b1212 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b1212 .OUTPUT_REG = 1'b0;
    defparam \RAM/MEM__D$b1212 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \RAM/MEM__D$b12c12  (.WCLK(\clk~O ), .RCLK(\clk~O ), .WCLKE(1'b1), 
            .WE(\RAM/n112 ), .RE(n107), .WDATA({\mem_wdata[19] }), .WADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RDATA({\RAM_rdata[19] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000010000000000000, INIT_1=256'h0000000000000300801002000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/bram/bram.v(12)
    defparam \RAM/MEM__D$b12c12 .READ_WIDTH = 1;
    defparam \RAM/MEM__D$b12c12 .WRITE_WIDTH = 1;
    defparam \RAM/MEM__D$b12c12 .WCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b12c12 .WCLKE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b12c12 .WE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b12c12 .RCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b12c12 .RE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b12c12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000010000000000000;
    defparam \RAM/MEM__D$b12c12 .INIT_1 = 256'h0000000000000300801002000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12c12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12c12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12c12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12c12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12c12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12c12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12c12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12c12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12c12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12c12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12c12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12c12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12c12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12c12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12c12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12c12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12c12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12c12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12c12 .OUTPUT_REG = 1'b0;
    defparam \RAM/MEM__D$b12c12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \RAM/MEM__D$b12d12  (.WCLK(\clk~O ), .RCLK(\clk~O ), .WCLKE(1'b1), 
            .WE(\RAM/n112 ), .RE(n107), .WDATA({\mem_wdata[20] }), .WADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RDATA({\RAM_rdata[20] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h032101400224204010030108004082111850401020C0400650500001E006B080, INIT_1=256'h00000000000064128B020428258018000060040040066C4AA880204C54400104, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/bram/bram.v(12)
    defparam \RAM/MEM__D$b12d12 .READ_WIDTH = 1;
    defparam \RAM/MEM__D$b12d12 .WRITE_WIDTH = 1;
    defparam \RAM/MEM__D$b12d12 .WCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b12d12 .WCLKE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b12d12 .WE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b12d12 .RCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b12d12 .RE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b12d12 .INIT_0 = 256'h032101400224204010030108004082111850401020C0400650500001E006B080;
    defparam \RAM/MEM__D$b12d12 .INIT_1 = 256'h00000000000064128B020428258018000060040040066C4AA880204C54400104;
    defparam \RAM/MEM__D$b12d12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12d12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12d12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12d12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12d12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12d12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12d12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12d12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12d12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12d12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12d12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12d12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12d12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12d12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12d12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12d12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12d12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12d12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12d12 .OUTPUT_REG = 1'b0;
    defparam \RAM/MEM__D$b12d12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \RAM/MEM__D$b12e12  (.WCLK(\clk~O ), .RCLK(\clk~O ), .WCLKE(1'b1), 
            .WE(\RAM/n112 ), .RE(n107), .WDATA({\mem_wdata[21] }), .WADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RDATA({\RAM_rdata[21] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h03210B80820500088002014009428A1150D1500020C20006B2000407A407A000, INIT_1=256'h0000000000006A1A6B405A18004010000260240240264848CC00204C76000804, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/bram/bram.v(12)
    defparam \RAM/MEM__D$b12e12 .READ_WIDTH = 1;
    defparam \RAM/MEM__D$b12e12 .WRITE_WIDTH = 1;
    defparam \RAM/MEM__D$b12e12 .WCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b12e12 .WCLKE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b12e12 .WE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b12e12 .RCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b12e12 .RE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b12e12 .INIT_0 = 256'h03210B80820500088002014009428A1150D1500020C20006B2000407A407A000;
    defparam \RAM/MEM__D$b12e12 .INIT_1 = 256'h0000000000006A1A6B405A18004010000260240240264848CC00204C76000804;
    defparam \RAM/MEM__D$b12e12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12e12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12e12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12e12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12e12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12e12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12e12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12e12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12e12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12e12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12e12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12e12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12e12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12e12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12e12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12e12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12e12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12e12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12e12 .OUTPUT_REG = 1'b0;
    defparam \RAM/MEM__D$b12e12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \RAM/MEM__D$b12f12  (.WCLK(\clk~O ), .RCLK(\clk~O ), .WCLKE(1'b1), 
            .WE(\RAM/n112 ), .RE(n107), .WDATA({\mem_wdata[22] }), .WADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RDATA({\RAM_rdata[22] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h07BB07A0532E01050086C7808D62CA1D51D1500134E00283E41A6EC5A0A6A001, INIT_1=256'h0000000000018F00E01358282504342083C83EA3C83CDD68F0047C6FD002A00F, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/bram/bram.v(12)
    defparam \RAM/MEM__D$b12f12 .READ_WIDTH = 1;
    defparam \RAM/MEM__D$b12f12 .WRITE_WIDTH = 1;
    defparam \RAM/MEM__D$b12f12 .WCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b12f12 .WCLKE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b12f12 .WE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b12f12 .RCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b12f12 .RE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b12f12 .INIT_0 = 256'h07BB07A0532E01050086C7808D62CA1D51D1500134E00283E41A6EC5A0A6A001;
    defparam \RAM/MEM__D$b12f12 .INIT_1 = 256'h0000000000018F00E01358282504342083C83EA3C83CDD68F0047C6FD002A00F;
    defparam \RAM/MEM__D$b12f12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12f12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12f12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12f12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12f12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12f12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12f12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12f12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12f12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12f12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12f12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12f12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12f12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12f12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12f12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12f12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12f12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12f12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12f12 .OUTPUT_REG = 1'b0;
    defparam \RAM/MEM__D$b12f12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \RAM/MEM__D$b12g1  (.WCLK(\clk~O ), .RCLK(\clk~O ), .WCLKE(1'b1), 
            .WE(\RAM/n112 ), .RE(n107), .WDATA({\mem_wdata[23] }), .WADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RDATA({\RAM_rdata[23] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h07FB4FA0E32F4329A18685D08D62CB1D55D5448330E28682A6980407B2A6E100, INIT_1=256'h000000000000002B17794219004C3630A2C82CA2EA2CD9D8FD0C784FDE86BA1F, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/bram/bram.v(12)
    defparam \RAM/MEM__D$b12g1 .READ_WIDTH = 1;
    defparam \RAM/MEM__D$b12g1 .WRITE_WIDTH = 1;
    defparam \RAM/MEM__D$b12g1 .WCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b12g1 .WCLKE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b12g1 .WE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b12g1 .RCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b12g1 .RE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$b12g1 .INIT_0 = 256'h07FB4FA0E32F4329A18685D08D62CB1D55D5448330E28682A6980407B2A6E100;
    defparam \RAM/MEM__D$b12g1 .INIT_1 = 256'h000000000000002B17794219004C3630A2C82CA2EA2CD9D8FD0C784FDE86BA1F;
    defparam \RAM/MEM__D$b12g1 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12g1 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12g1 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12g1 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12g1 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12g1 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12g1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12g1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12g1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12g1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12g1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12g1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12g1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12g1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12g1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12g1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12g1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12g1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$b12g1 .OUTPUT_REG = 1'b0;
    defparam \RAM/MEM__D$b12g1 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \RAM/MEM__D$1212  (.WCLK(\clk~O ), .RCLK(\clk~O ), .WCLKE(1'b1), 
            .WE(\RAM/n108 ), .RE(n107), .WDATA({\mem_wdata[9] }), .WADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RDATA({\RAM_rdata[9] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h1FBB85F8431F2040900F8DC83EFDF7EFBE7EF68018F2401FFE40C38FE047BC90, INIT_1=256'h00000000000000142A9CCBB23A81FC6187F87F87F87FF776AC80F8FF7A400907, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/bram/bram.v(12)
    defparam \RAM/MEM__D$1212 .READ_WIDTH = 1;
    defparam \RAM/MEM__D$1212 .WRITE_WIDTH = 1;
    defparam \RAM/MEM__D$1212 .WCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$1212 .WCLKE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$1212 .WE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$1212 .RCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$1212 .RE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$1212 .INIT_0 = 256'h1FBB85F8431F2040900F8DC83EFDF7EFBE7EF68018F2401FFE40C38FE047BC90;
    defparam \RAM/MEM__D$1212 .INIT_1 = 256'h00000000000000142A9CCBB23A81FC6187F87F87F87FF776AC80F8FF7A400907;
    defparam \RAM/MEM__D$1212 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$1212 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$1212 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$1212 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$1212 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$1212 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$1212 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$1212 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$1212 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$1212 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$1212 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$1212 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$1212 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$1212 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$1212 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$1212 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$1212 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$1212 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$1212 .OUTPUT_REG = 1'b0;
    defparam \RAM/MEM__D$1212 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \RAM/MEM__D$12c12  (.WCLK(\clk~O ), .RCLK(\clk~O ), .WCLKE(1'b1), 
            .WE(\RAM/n108 ), .RE(n107), .WDATA({\mem_wdata[11] }), .WADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RDATA({\RAM_rdata[11] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h00050000001100003010004001020800001008802002000000C0000400000180, INIT_1=256'h0000000000009B94080A808445001000000000000000400BC400000006000304, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/bram/bram.v(12)
    defparam \RAM/MEM__D$12c12 .READ_WIDTH = 1;
    defparam \RAM/MEM__D$12c12 .WRITE_WIDTH = 1;
    defparam \RAM/MEM__D$12c12 .WCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$12c12 .WCLKE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$12c12 .WE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$12c12 .RCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$12c12 .RE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$12c12 .INIT_0 = 256'h00050000001100003010004001020800001008802002000000C0000400000180;
    defparam \RAM/MEM__D$12c12 .INIT_1 = 256'h0000000000009B94080A808445001000000000000000400BC400000006000304;
    defparam \RAM/MEM__D$12c12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12c12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12c12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12c12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12c12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12c12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12c12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12c12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12c12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12c12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12c12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12c12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12c12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12c12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12c12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12c12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12c12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12c12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12c12 .OUTPUT_REG = 1'b0;
    defparam \RAM/MEM__D$12c12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \RAM/MEM__D$12d12  (.WCLK(\clk~O ), .RCLK(\clk~O ), .WCLKE(1'b1), 
            .WE(\RAM/n108 ), .RE(n107), .WDATA({\mem_wdata[12] }), .WADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RDATA({\RAM_rdata[12] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0004010000100000001000000000001010104800000000055010000400000002, INIT_1=256'h000000000000E0140A88840A6000800000400400400408000000800C20000004, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/bram/bram.v(12)
    defparam \RAM/MEM__D$12d12 .READ_WIDTH = 1;
    defparam \RAM/MEM__D$12d12 .WRITE_WIDTH = 1;
    defparam \RAM/MEM__D$12d12 .WCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$12d12 .WCLKE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$12d12 .WE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$12d12 .RCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$12d12 .RE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$12d12 .INIT_0 = 256'h0004010000100000001000000000001010104800000000055010000400000002;
    defparam \RAM/MEM__D$12d12 .INIT_1 = 256'h000000000000E0140A88840A6000800000400400400408000000800C20000004;
    defparam \RAM/MEM__D$12d12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12d12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12d12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12d12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12d12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12d12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12d12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12d12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12d12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12d12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12d12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12d12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12d12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12d12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12d12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12d12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12d12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12d12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12d12 .OUTPUT_REG = 1'b0;
    defparam \RAM/MEM__D$12d12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \RAM/MEM__D$12e12  (.WCLK(\clk~O ), .RCLK(\clk~O ), .WCLKE(1'b1), 
            .WE(\RAM/n108 ), .RE(n107), .WDATA({\mem_wdata[13] }), .WADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RDATA({\RAM_rdata[13] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h069305A0410D6301B18685D8AD2A695DC485648330A2C60006D1040400000182, INIT_1=256'h000000000000EE100A09800B354C3420868868868868D15BFD8C680B4EC62B1A, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/bram/bram.v(12)
    defparam \RAM/MEM__D$12e12 .READ_WIDTH = 1;
    defparam \RAM/MEM__D$12e12 .WRITE_WIDTH = 1;
    defparam \RAM/MEM__D$12e12 .WCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$12e12 .WCLKE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$12e12 .WE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$12e12 .RCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$12e12 .RE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$12e12 .INIT_0 = 256'h069305A0410D6301B18685D8AD2A695DC485648330A2C60006D1040400000182;
    defparam \RAM/MEM__D$12e12 .INIT_1 = 256'h000000000000EE100A09800B354C3420868868868868D15BFD8C680B4EC62B1A;
    defparam \RAM/MEM__D$12e12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12e12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12e12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12e12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12e12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12e12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12e12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12e12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12e12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12e12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12e12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12e12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12e12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12e12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12e12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12e12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12e12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12e12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12e12 .OUTPUT_REG = 1'b0;
    defparam \RAM/MEM__D$12e12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \RAM/MEM__D$12f12  (.WCLK(\clk~O ), .RCLK(\clk~O ), .WCLKE(1'b1), 
            .WE(\RAM/n108 ), .RE(n107), .WDATA({\mem_wdata[14] }), .WADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RDATA({\RAM_rdata[14] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0800010000100000000808000000001000004000200000000010000520048000, INIT_1=256'h0000000000010A2414898D8A2000404100100100100102000000808C00000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/bram/bram.v(12)
    defparam \RAM/MEM__D$12f12 .READ_WIDTH = 1;
    defparam \RAM/MEM__D$12f12 .WRITE_WIDTH = 1;
    defparam \RAM/MEM__D$12f12 .WCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$12f12 .WCLKE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$12f12 .WE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$12f12 .RCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$12f12 .RE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$12f12 .INIT_0 = 256'h0800010000100000000808000000001000004000200000000010000520048000;
    defparam \RAM/MEM__D$12f12 .INIT_1 = 256'h0000000000010A2414898D8A2000404100100100100102000000808C00000000;
    defparam \RAM/MEM__D$12f12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12f12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12f12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12f12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12f12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12f12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12f12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12f12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12f12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12f12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12f12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12f12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12f12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12f12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12f12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12f12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12f12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12f12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12f12 .OUTPUT_REG = 1'b0;
    defparam \RAM/MEM__D$12f12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \RAM/MEM__D$12g1  (.WCLK(\clk~O ), .RCLK(\clk~O ), .WCLKE(1'b1), 
            .WE(\RAM/n108 ), .RE(n107), .WDATA({\mem_wdata[15] }), .WADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RDATA({\RAM_rdata[15] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'hB9045355149008A404195802692A294444856C28040810A9F019A55452A90008, INIT_1=256'h000000000000000122BF83459562CACB2D12D12D12D122200020958830108040, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/bram/bram.v(12)
    defparam \RAM/MEM__D$12g1 .READ_WIDTH = 1;
    defparam \RAM/MEM__D$12g1 .WRITE_WIDTH = 1;
    defparam \RAM/MEM__D$12g1 .WCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$12g1 .WCLKE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$12g1 .WE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$12g1 .RCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$12g1 .RE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$12g1 .INIT_0 = 256'hB9045355149008A404195802692A294444856C28040810A9F019A55452A90008;
    defparam \RAM/MEM__D$12g1 .INIT_1 = 256'h000000000000000122BF83459562CACB2D12D12D12D122200020958830108040;
    defparam \RAM/MEM__D$12g1 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12g1 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12g1 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12g1 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12g1 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12g1 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12g1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12g1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12g1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12g1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12g1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12g1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12g1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12g1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12g1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12g1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12g1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12g1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$12g1 .OUTPUT_REG = 1'b0;
    defparam \RAM/MEM__D$12g1 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \RAM/MEM__D$212  (.WCLK(\clk~O ), .RCLK(\clk~O ), .WCLKE(1'b1), 
            .WE(\RAM/n104 ), .RE(n107), .WDATA({\mem_wdata[1] }), .WADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RDATA({\RAM_rdata[1] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_1=256'h0000000000011D8F21F1D3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/bram/bram.v(12)
    defparam \RAM/MEM__D$212 .READ_WIDTH = 1;
    defparam \RAM/MEM__D$212 .WRITE_WIDTH = 1;
    defparam \RAM/MEM__D$212 .WCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$212 .WCLKE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$212 .WE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$212 .RCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$212 .RE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$212 .INIT_0 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \RAM/MEM__D$212 .INIT_1 = 256'h0000000000011D8F21F1D3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \RAM/MEM__D$212 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$212 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$212 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$212 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$212 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$212 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$212 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$212 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$212 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$212 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$212 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$212 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$212 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$212 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$212 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$212 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$212 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$212 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$212 .OUTPUT_REG = 1'b0;
    defparam \RAM/MEM__D$212 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \RAM/MEM__D$2c12  (.WCLK(\clk~O ), .RCLK(\clk~O ), .WCLKE(1'b1), 
            .WE(\RAM/n104 ), .RE(n107), .WDATA({\mem_wdata[3] }), .WADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RDATA({\RAM_rdata[3] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0040000020000000000002000000000001000000000000000010000000004000, INIT_1=256'h0000000000009381002006000000001040040040040000800000000080000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/bram/bram.v(12)
    defparam \RAM/MEM__D$2c12 .READ_WIDTH = 1;
    defparam \RAM/MEM__D$2c12 .WRITE_WIDTH = 1;
    defparam \RAM/MEM__D$2c12 .WCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$2c12 .WCLKE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$2c12 .WE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$2c12 .RCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$2c12 .RE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$2c12 .INIT_0 = 256'h0040000020000000000002000000000001000000000000000010000000004000;
    defparam \RAM/MEM__D$2c12 .INIT_1 = 256'h0000000000009381002006000000001040040040040000800000000080000000;
    defparam \RAM/MEM__D$2c12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2c12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2c12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2c12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2c12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2c12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2c12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2c12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2c12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2c12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2c12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2c12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2c12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2c12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2c12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2c12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2c12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2c12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2c12 .OUTPUT_REG = 1'b0;
    defparam \RAM/MEM__D$2c12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \RAM/MEM__D$2d12  (.WCLK(\clk~O ), .RCLK(\clk~O ), .WCLKE(1'b1), 
            .WE(\RAM/n104 ), .RE(n107), .WDATA({\mem_wdata[4] }), .WADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RDATA({\RAM_rdata[4] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h7108B95B8E6294DA4A61302552D596A2BA6AD354CB55297FF926DBBA4DD91257, INIT_1=256'h000000000000E83A054A941A2A93098619219219219224240253137C312954A1, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/bram/bram.v(12)
    defparam \RAM/MEM__D$2d12 .READ_WIDTH = 1;
    defparam \RAM/MEM__D$2d12 .WRITE_WIDTH = 1;
    defparam \RAM/MEM__D$2d12 .WCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$2d12 .WCLKE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$2d12 .WE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$2d12 .RCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$2d12 .RE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$2d12 .INIT_0 = 256'h7108B95B8E6294DA4A61302552D596A2BA6AD354CB55297FF926DBBA4DD91257;
    defparam \RAM/MEM__D$2d12 .INIT_1 = 256'h000000000000E83A054A941A2A93098619219219219224240253137C312954A1;
    defparam \RAM/MEM__D$2d12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2d12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2d12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2d12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2d12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2d12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2d12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2d12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2d12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2d12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2d12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2d12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2d12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2d12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2d12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2d12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2d12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2d12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2d12 .OUTPUT_REG = 1'b0;
    defparam \RAM/MEM__D$2d12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \RAM/MEM__D$2e12  (.WCLK(\clk~O ), .RCLK(\clk~O ), .WCLKE(1'b1), 
            .WE(\RAM/n104 ), .RE(n107), .WDATA({\mem_wdata[5] }), .WADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RDATA({\RAM_rdata[5] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h8265428432956824B412435A1BD79EB3F3B39AB824CAD082A2D964CC92626DAB, INIT_1=256'h000000000000EA2F1DE997E4E560921862462462462448CBFDA0A454C6D08B44, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/bram/bram.v(12)
    defparam \RAM/MEM__D$2e12 .READ_WIDTH = 1;
    defparam \RAM/MEM__D$2e12 .WRITE_WIDTH = 1;
    defparam \RAM/MEM__D$2e12 .WCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$2e12 .WCLKE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$2e12 .WE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$2e12 .RCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$2e12 .RE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$2e12 .INIT_0 = 256'h8265428432956824B412435A1BD79EB3F3B39AB824CAD082A2D964CC92626DAB;
    defparam \RAM/MEM__D$2e12 .INIT_1 = 256'h000000000000EA2F1DE997E4E560921862462462462448CBFDA0A454C6D08B44;
    defparam \RAM/MEM__D$2e12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2e12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2e12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2e12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2e12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2e12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2e12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2e12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2e12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2e12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2e12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2e12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2e12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2e12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2e12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2e12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2e12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2e12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2e12 .OUTPUT_REG = 1'b0;
    defparam \RAM/MEM__D$2e12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \RAM/MEM__D$2f12  (.WCLK(\clk~O ), .RCLK(\clk~O ), .WCLKE(1'b1), 
            .WE(\RAM/n104 ), .RE(n107), .WDATA({\mem_wdata[6] }), .WADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RDATA({\RAM_rdata[6] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h8064400430900824041042020000001081100838240810800018204412204028, INIT_1=256'h0000000000010E140A8925E4C020821860460460460408800020840080108044, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/bram/bram.v(12)
    defparam \RAM/MEM__D$2f12 .READ_WIDTH = 1;
    defparam \RAM/MEM__D$2f12 .WRITE_WIDTH = 1;
    defparam \RAM/MEM__D$2f12 .WCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$2f12 .WCLKE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$2f12 .WE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$2f12 .RCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$2f12 .RE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$2f12 .INIT_0 = 256'h8064400430900824041042020000001081100838240810800018204412204028;
    defparam \RAM/MEM__D$2f12 .INIT_1 = 256'h0000000000010E140A8925E4C020821860460460460408800020840080108044;
    defparam \RAM/MEM__D$2f12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2f12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2f12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2f12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2f12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2f12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2f12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2f12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2f12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2f12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2f12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2f12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2f12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2f12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2f12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2f12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2f12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2f12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2f12 .OUTPUT_REG = 1'b0;
    defparam \RAM/MEM__D$2f12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \RAM/MEM__D$2g1  (.WCLK(\clk~O ), .RCLK(\clk~O ), .WCLKE(1'b1), 
            .WE(\RAM/n104 ), .RE(n107), .WDATA({\mem_wdata[7] }), .WADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RADDR({\mem_addr[13] , 
            \mem_addr[12] , \mem_addr[11] , \mem_addr[10] , \mem_addr[9] , 
            \mem_addr[8] , \mem_addr[7] , \mem_addr[6] , \mem_addr[5] , 
            \mem_addr[4] , \mem_addr[3] , \mem_addr[2] }), .RDATA({\RAM_rdata[7] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'hDDAEEC3EDBCA0176009DEC8032B555A6A62AB601366C02D4F80CF1EEFB75B40D, INIT_1=256'h0000000000000026371EF8364A85EF6DB4AB4AB4AB4AB5340004DECD3802D00D, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/bram/bram.v(12)
    defparam \RAM/MEM__D$2g1 .READ_WIDTH = 1;
    defparam \RAM/MEM__D$2g1 .WRITE_WIDTH = 1;
    defparam \RAM/MEM__D$2g1 .WCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$2g1 .WCLKE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$2g1 .WE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$2g1 .RCLK_POLARITY = 1'b1;
    defparam \RAM/MEM__D$2g1 .RE_POLARITY = 1'b1;
    defparam \RAM/MEM__D$2g1 .INIT_0 = 256'hDDAEEC3EDBCA0176009DEC8032B555A6A62AB601366C02D4F80CF1EEFB75B40D;
    defparam \RAM/MEM__D$2g1 .INIT_1 = 256'h0000000000000026371EF8364A85EF6DB4AB4AB4AB4AB5340004DECD3802D00D;
    defparam \RAM/MEM__D$2g1 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2g1 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2g1 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2g1 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2g1 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2g1 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2g1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2g1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2g1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2g1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2g1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2g1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2g1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2g1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2g1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2g1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2g1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2g1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \RAM/MEM__D$2g1 .OUTPUT_REG = 1'b0;
    defparam \RAM/MEM__D$2g1 .WRITE_MODE = "READ_FIRST";
    EFX_LUT4 LUT__2369 (.I0(\mem_wdata[0] ), .I1(\CPU/instr[20] ), .I2(\CPU/instr[4]~FF_frt_1_q ), 
            .I3(\CPU/instr[2]~FF_frt_0_q ), .O(n1587)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__2369.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__2370 (.I0(\CPU/instr[4] ), .I1(\CPU/instr[8] ), .I2(\CPU/instr[21] ), 
            .I3(\CPU/instr[3] ), .O(n787)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044 */ ;
    defparam LUT__2370.LUTMASK = 16'hf044;
    EFX_LUT4 LUT__2371 (.I0(\CPU/aluShamt[0] ), .I1(\CPU/aluShamt[1] ), 
            .I2(\CPU/aluShamt[2] ), .O(n1590)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__2371.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__2372 (.I0(\CPU/aluShamt[3] ), .I1(n1590), .O(n1591)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2372.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2373 (.I0(\CPU/aluShamt[4] ), .I1(n1591), .O(n1592)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2373.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2374 (.I0(n1587), .I1(n1592), .I2(\CPU/aluShamt[0] ), 
            .O(\CPU/n1034 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__2374.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__2375 (.I0(\CPU/instr[2] ), .I1(\CPU/instr[3] ), .I2(\CPU/instr[6] ), 
            .I3(\CPU/instr[4] ), .O(n1593)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__2375.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__2376 (.I0(\CPU/instr[13] ), .I1(\CPU/instr[12] ), .O(n1594)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2376.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2377 (.I0(n1593), .I1(n1594), .O(n1595)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2377.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2378 (.I0(\CPU/state[2] ), .I1(n1595), .I2(n1592), .O(ceg_net77)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2378.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2379 (.I0(\CPU/instr[2] ), .I1(\CPU/instr[3] ), .O(n1596)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__2379.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__2380 (.I0(\CPU/instr[4] ), .I1(n1594), .I2(\CPU/instr[6] ), 
            .I3(n1596), .O(n1597)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__2380.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__2381 (.I0(\CPU/state[0] ), .I1(n1592), .I2(\CPU/state[3] ), 
            .O(n1598)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__2381.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__2382 (.I0(n1597), .I1(\CPU/state[2] ), .I2(n1598), .O(\CPU/n2185 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__2382.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__2383 (.I0(\CPU/instr[20] ), .I1(\CPU/instr[7] ), .I2(\CPU/instr[5] ), 
            .O(n793)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__2383.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__2384 (.I0(\CPU/instr[4] ), .I1(\CPU/instr[5] ), .I2(\CPU/instr[6] ), 
            .I3(n1596), .O(n1599)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__2384.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__2385 (.I0(n580), .I1(\CPU/PC[17] ), .I2(\CPU/state[0] ), 
            .I3(\CPU/state[1] ), .O(n1600)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca */ ;
    defparam LUT__2385.LUTMASK = 16'hccca;
    EFX_LUT4 LUT__2386 (.I0(n578), .I1(\CPU/PC[18] ), .I2(\CPU/state[0] ), 
            .I3(\CPU/state[1] ), .O(n1601)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca */ ;
    defparam LUT__2386.LUTMASK = 16'hccca;
    EFX_LUT4 LUT__2387 (.I0(n1600), .I1(n1601), .O(n1602)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2387.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2388 (.I0(n576), .I1(\CPU/PC[19] ), .I2(\CPU/state[0] ), 
            .I3(\CPU/state[1] ), .O(n1603)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca */ ;
    defparam LUT__2388.LUTMASK = 16'hccca;
    EFX_LUT4 LUT__2389 (.I0(n569), .I1(n572), .I2(n574), .O(n1604)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__2389.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__2390 (.I0(\CPU/PC[20] ), .I1(\CPU/PC[21] ), .I2(\CPU/PC[23] ), 
            .O(n1605)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__2390.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__2391 (.I0(\CPU/state[0] ), .I1(\CPU/state[1] ), .O(n1606)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__2391.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__2392 (.I0(n570), .I1(\CPU/PC[22] ), .I2(\CPU/state[0] ), 
            .I3(\CPU/state[1] ), .O(n1607)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3335 */ ;
    defparam LUT__2392.LUTMASK = 16'h3335;
    EFX_LUT4 LUT__2393 (.I0(n1605), .I1(n1604), .I2(n1607), .I3(n1606), 
            .O(n1608)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__2393.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__2394 (.I0(n1602), .I1(n1603), .I2(n1608), .O(n1609)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__2394.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__2395 (.I0(n1599), .I1(\CPU/state[2] ), .I2(\CPU/state[0] ), 
            .I3(n1609), .O(n107)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f8 */ ;
    defparam LUT__2395.LUTMASK = 16'h00f8;
    EFX_LUT4 LUT__2396 (.I0(\CPU/PC[2] ), .I1(n610), .I2(n1606), .O(\mem_addr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__2396.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__2397 (.I0(\CPU/PC[3] ), .I1(n608), .I2(n1606), .O(\mem_addr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__2397.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__2398 (.I0(\CPU/PC[4] ), .I1(n606), .I2(n1606), .O(\mem_addr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__2398.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__2399 (.I0(\CPU/PC[5] ), .I1(n604), .I2(n1606), .O(\mem_addr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__2399.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__2400 (.I0(\CPU/PC[6] ), .I1(n602), .I2(n1606), .O(\mem_addr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__2400.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__2401 (.I0(\CPU/PC[7] ), .I1(n600), .I2(n1606), .O(\mem_addr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__2401.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__2402 (.I0(\CPU/PC[8] ), .I1(n598), .I2(n1606), .O(\mem_addr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__2402.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__2403 (.I0(\CPU/PC[9] ), .I1(n596), .I2(n1606), .O(\mem_addr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__2403.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__2404 (.I0(\CPU/PC[10] ), .I1(n594), .I2(n1606), .O(\mem_addr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__2404.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__2405 (.I0(\CPU/PC[11] ), .I1(n592), .I2(n1606), .O(\mem_addr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__2405.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__2406 (.I0(\CPU/PC[12] ), .I1(n590), .I2(n1606), .O(\mem_addr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__2406.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__2407 (.I0(\CPU/PC[13] ), .I1(n588), .I2(n1606), .O(\mem_addr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__2407.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__2408 (.I0(\CPU/rs2[8] ), .I1(\mem_wdata[0] ), .I2(n12), 
            .O(\mem_wdata[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__2408.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__2409 (.I0(n12), .I1(n612), .O(n1610)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__2409.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__2410 (.I0(\mem_wdata[8] ), .I1(\CPU/rs2[24] ), .I2(n1610), 
            .O(\mem_wdata[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__2410.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__2411 (.I0(\CPU/instr[12] ), .I1(\CPU/instr[13] ), .O(n1611)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__2411.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__2412 (.I0(\CPU/instr[4] ), .I1(\CPU/instr[6] ), .I2(\CPU/instr[2]~FF_frt_0_q ), 
            .I3(\CPU/state[2] ), .O(n1612)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__2412.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__2413 (.I0(n582), .I1(\CPU/PC[16] ), .I2(\CPU/state[0] ), 
            .I3(\CPU/state[1] ), .O(n1613)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3335 */ ;
    defparam LUT__2413.LUTMASK = 16'h3335;
    EFX_LUT4 LUT__2414 (.I0(n1603), .I1(n1601), .I2(n1613), .O(n1614)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__2414.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__2415 (.I0(n1600), .I1(n1612), .I2(n1614), .O(n1615)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__2415.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__2416 (.I0(\CPU/PC[14] ), .I1(\CPU/PC[15] ), .I2(\CPU/PC[22] ), 
            .O(n1616)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__2416.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__2417 (.I0(n570), .I1(n584), .I2(n586), .O(n1617)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__2417.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__2418 (.I0(n1604), .I1(n1617), .I2(n1616), .I3(n1606), 
            .O(n1618)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f */ ;
    defparam LUT__2418.LUTMASK = 16'h770f;
    EFX_LUT4 LUT__2419 (.I0(n1606), .I1(n1605), .I2(n1618), .I3(n1615), 
            .O(n1619)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__2419.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__2420 (.I0(n612), .I1(\CPU/instr[13] ), .I2(n1619), .O(n1620)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__2420.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__2421 (.I0(n12), .I1(n1611), .I2(n1620), .O(\RAM/n116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__2421.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__2422 (.I0(resetn), .I1(\CPU/state[1] ), .O(\CPU/n3447 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2422.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2423 (.I0(n1601), .I1(n1603), .I2(n1600), .I3(n1613), 
            .O(n1621)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__2423.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__2424 (.I0(n1608), .I1(n1621), .O(n1622)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2424.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2425 (.I0(n1603), .I1(n1602), .I2(n1608), .I3(\RAM_rdata[15] ), 
            .O(n1623)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__2425.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__2426 (.I0(n1622), .I1(\mult_dout[15] ), .I2(n1623), 
            .O(\mem_rdata[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8 */ ;
    defparam LUT__2426.LUTMASK = 16'hf8f8;
    EFX_LUT4 LUT__2427 (.I0(n1622), .I1(\mult_dout[16] ), .I2(n1609), 
            .I3(\RAM_rdata[16] ), .O(\mem_rdata[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f88 */ ;
    defparam LUT__2427.LUTMASK = 16'h8f88;
    EFX_LUT4 LUT__2428 (.I0(n1622), .I1(\mult_dout[17] ), .I2(n1609), 
            .I3(\RAM_rdata[17] ), .O(\mem_rdata[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f88 */ ;
    defparam LUT__2428.LUTMASK = 16'h8f88;
    EFX_LUT4 LUT__2429 (.I0(n1622), .I1(\mult_dout[18] ), .I2(n1609), 
            .I3(\RAM_rdata[18] ), .O(\mem_rdata[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f88 */ ;
    defparam LUT__2429.LUTMASK = 16'h8f88;
    EFX_LUT4 LUT__2430 (.I0(n1608), .I1(n1621), .I2(\mult_dout[19] ), 
            .O(n1624)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__2430.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__2431 (.I0(n1609), .I1(\RAM_rdata[19] ), .I2(n1624), 
            .O(\mem_rdata[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__2431.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__2432 (.I0(n1608), .I1(n1621), .I2(\mult_dout[23] ), 
            .O(n1625)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__2432.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__2433 (.I0(n12), .I1(n1611), .I2(n612), .O(n1626)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__2433.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__2434 (.I0(\RAM_rdata[23] ), .I1(n1609), .I2(n1625), 
            .I3(n1626), .O(n1627)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__2434.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__2435 (.I0(n12), .I1(n1611), .I2(n612), .O(n1628)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__2435.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__2436 (.I0(\mult_dout[15] ), .I1(n1621), .I2(n1608), 
            .I3(n1628), .O(n1629)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00 */ ;
    defparam LUT__2436.LUTMASK = 16'h7f00;
    EFX_LUT4 LUT__2437 (.I0(n1603), .I1(n1602), .I2(n1608), .I3(\RAM_rdata[31] ), 
            .O(n1630)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__2437.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__2438 (.I0(n12), .I1(n1611), .I2(n612), .O(n1631)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__2438.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__2439 (.I0(\mult_dout[31] ), .I1(n1621), .I2(n1608), 
            .I3(n1631), .O(n1632)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00 */ ;
    defparam LUT__2439.LUTMASK = 16'h7f00;
    EFX_LUT4 LUT__2440 (.I0(n1630), .I1(n1632), .I2(n1623), .I3(n1629), 
            .O(n1633)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__2440.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__2441 (.I0(n1603), .I1(n1602), .I2(n1608), .I3(\RAM_rdata[7] ), 
            .O(n1634)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__2441.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__2442 (.I0(\uart_dout[7] ), .I1(\mult_dout[7] ), .I2(n1600), 
            .O(n1635)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__2442.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__2443 (.I0(n1635), .I1(n1614), .I2(n1608), .O(n1636)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__2443.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__2444 (.I0(n1610), .I1(n1611), .O(n1637)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2444.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2445 (.I0(\CPU/instr[14] ), .I1(n1599), .O(n1638)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2445.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2446 (.I0(n1636), .I1(n1634), .I2(n1637), .I3(n1638), 
            .O(n1639)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__2446.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__2447 (.I0(n1627), .I1(\CPU/instr[13] ), .I2(n1633), 
            .I3(n1639), .O(n1640)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__2447.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__2448 (.I0(n703), .I1(n705), .I2(n707), .I3(n717), 
            .O(n1641)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2448.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2449 (.I0(n709), .I1(n711), .I2(n713), .I3(n715), 
            .O(n1642)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2449.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2450 (.I0(n693), .I1(n695), .I2(n697), .I3(n699), 
            .O(n1643)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2450.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2451 (.I0(n6), .I1(n689), .I2(n691), .I3(n701), .O(n1644)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2451.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2452 (.I0(n1641), .I1(n1642), .I2(n1643), .I3(n1644), 
            .O(n1645)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2452.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2453 (.I0(\CPU/instr[5] ), .I1(\CPU/instr[30] ), .O(n1646)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2453.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2454 (.I0(n748), .I1(n687), .I2(n1645), .I3(n1646), 
            .O(n1647)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc355 */ ;
    defparam LUT__2454.LUTMASK = 16'hc355;
    EFX_LUT4 LUT__2455 (.I0(\CPU/rs2[16] ), .I1(\CPU/instr[31] ), .I2(\CPU/instr[4]~FF_frt_1_q ), 
            .I3(\CPU/instr[2]~FF_frt_0_q ), .O(n1555)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__2455.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__2456 (.I0(n1647), .I1(n1555), .I2(\CPU/rs1[16] ), .I3(\CPU/instr[14] ), 
            .O(n1648)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3c55 */ ;
    defparam LUT__2456.LUTMASK = 16'h3c55;
    EFX_LUT4 LUT__2457 (.I0(\CPU/instr[13] ), .I1(\CPU/instr[14] ), .O(n1649)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2457.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2458 (.I0(n1555), .I1(\CPU/instr[12] ), .I2(\CPU/rs1[16] ), 
            .I3(n1649), .O(n1650)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb200 */ ;
    defparam LUT__2458.LUTMASK = 16'hb200;
    EFX_LUT4 LUT__2459 (.I0(\CPU/aluReg[16] ), .I1(n1594), .I2(n1650), 
            .O(n1651)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__2459.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__2460 (.I0(n1611), .I1(n1648), .I2(n1651), .I3(n1593), 
            .O(n1652)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__2460.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__2461 (.I0(n1599), .I1(\CPU/instr[13] ), .O(n1653)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2461.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2462 (.I0(\CPU/instr[3] ), .I1(\CPU/instr[2] ), .O(n1654)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2462.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2463 (.I0(\CPU/instr[6] ), .I1(\CPU/instr[4] ), .O(n1655)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2463.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2464 (.I0(\CPU/instr[5] ), .I1(n1654), .I2(n1655), .O(n1656)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__2464.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__2465 (.I0(n1656), .I1(n627), .I2(\mem_rdata[16] ), .I3(n1653), 
            .O(n1657)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2465.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2466 (.I0(\CPU/PC[2] ), .I1(\CPU/PC[3] ), .I2(\CPU/PC[4] ), 
            .I3(\CPU/PC[5] ), .O(n1658)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2466.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2467 (.I0(\CPU/PC[10] ), .I1(\CPU/PC[11] ), .I2(\CPU/PC[12] ), 
            .I3(\CPU/PC[13] ), .O(n1659)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2467.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2468 (.I0(\CPU/PC[6] ), .I1(\CPU/PC[7] ), .I2(\CPU/PC[8] ), 
            .I3(\CPU/PC[9] ), .O(n1660)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2468.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2469 (.I0(n1658), .I1(n1659), .I2(n1660), .O(n1661)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__2469.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__2470 (.I0(n1661), .I1(\CPU/PC[14] ), .I2(\CPU/PC[15] ), 
            .I3(\CPU/PC[16] ), .O(n1662)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__2470.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__2471 (.I0(\CPU/instr[4] ), .I1(\CPU/instr[5] ), .I2(\CPU/instr[6] ), 
            .O(n1663)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__2471.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__2472 (.I0(\CPU/instr[2] ), .I1(n1663), .I2(\CPU/instr[3] ), 
            .O(n1664)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__2472.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__2473 (.I0(\CPU/instr[2]~FF_frt_0_q ), .I1(\CPU/instr[4] ), 
            .I2(\CPU/instr[6] ), .O(n1665)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__2473.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__2474 (.I0(n1655), .I1(n1654), .I2(\CPU/instr[5] ), .O(n1666)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__2474.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__2475 (.I0(\CPU/instr[16] ), .I1(n1666), .I2(n1665), 
            .I3(\CPU/cycles[16] ), .O(n1667)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2475.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2476 (.I0(n1664), .I1(n1662), .I2(n1667), .O(n1668)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__2476.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__2477 (.I0(n1640), .I1(n1652), .I2(n1657), .I3(n1668), 
            .O(\CPU/writeBackData[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hefff */ ;
    defparam LUT__2477.LUTMASK = 16'hefff;
    EFX_LUT4 LUT__2478 (.I0(n1645), .I1(n687), .I2(n685), .I3(n1646), 
            .O(n1669)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8700 */ ;
    defparam LUT__2478.LUTMASK = 16'h8700;
    EFX_LUT4 LUT__2479 (.I0(\CPU/instr[12] ), .I1(\CPU/instr[13] ), .I2(\CPU/instr[14] ), 
            .O(n1670)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__2479.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__2480 (.I0(n746), .I1(n1646), .I2(n1669), .I3(n1670), 
            .O(n1671)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__2480.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__2481 (.I0(n1594), .I1(\CPU/aluReg[17] ), .O(n1672)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2481.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2482 (.I0(\CPU/instr[12] ), .I1(\CPU/instr[14] ), .O(n1673)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2482.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2483 (.I0(n1588), .I1(n1589), .O(n1674)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2483.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2484 (.I0(\CPU/instr[31] ), .I1(\CPU/rs2[17] ), .I2(\CPU/instr[4]~FF_frt_1_frt_2_q ), 
            .O(n1553)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__2484.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__2485 (.I0(n1649), .I1(n1673), .I2(n1553), .I3(\CPU/rs1[17] ), 
            .O(n1675)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h533f */ ;
    defparam LUT__2485.LUTMASK = 16'h533f;
    EFX_LUT4 LUT__2486 (.I0(n1672), .I1(n1671), .I2(n1675), .I3(n1593), 
            .O(n1676)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__2486.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__2487 (.I0(\CPU/PC[14] ), .I1(\CPU/PC[15] ), .I2(\CPU/PC[16] ), 
            .O(n1677)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__2487.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__2488 (.I0(n1661), .I1(n1677), .I2(n1664), .I3(\CPU/PC[17] ), 
            .O(n1678)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0708 */ ;
    defparam LUT__2488.LUTMASK = 16'h0708;
    EFX_LUT4 LUT__2489 (.I0(n1656), .I1(n625), .I2(n1665), .I3(\CPU/cycles[17] ), 
            .O(n1679)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2489.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2490 (.I0(\CPU/instr[17] ), .I1(n1666), .I2(n1678), 
            .I3(n1679), .O(n1680)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__2490.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__2491 (.I0(n1653), .I1(\mem_rdata[17] ), .I2(n1680), 
            .O(n1681)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2491.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2492 (.I0(n1640), .I1(n1676), .I2(n1681), .O(\CPU/writeBackData[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hefef */ ;
    defparam LUT__2492.LUTMASK = 16'hefef;
    EFX_LUT4 LUT__2493 (.I0(n685), .I1(n687), .O(n1682)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2493.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2494 (.I0(n1645), .I1(n1682), .I2(n683), .I3(n1646), 
            .O(n1683)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8700 */ ;
    defparam LUT__2494.LUTMASK = 16'h8700;
    EFX_LUT4 LUT__2495 (.I0(n744), .I1(n1646), .I2(n1670), .O(n1684)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__2495.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__2496 (.I0(\CPU/rs2[18] ), .I1(\CPU/instr[31] ), .I2(\CPU/instr[4]~FF_frt_1_q ), 
            .I3(\CPU/instr[2]~FF_frt_0_q ), .O(n1551)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__2496.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__2497 (.I0(\CPU/instr[13] ), .I1(\CPU/instr[12] ), .I2(n1551), 
            .I3(\CPU/rs1[18] ), .O(n1685)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ccf */ ;
    defparam LUT__2497.LUTMASK = 16'h5ccf;
    EFX_LUT4 LUT__2498 (.I0(n1594), .I1(\CPU/aluReg[18] ), .I2(n1685), 
            .I3(\CPU/instr[14] ), .O(n1686)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077 */ ;
    defparam LUT__2498.LUTMASK = 16'h7077;
    EFX_LUT4 LUT__2499 (.I0(n1683), .I1(n1684), .I2(n1686), .I3(n1593), 
            .O(n1687)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__2499.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__2500 (.I0(\CPU/PC[14] ), .I1(\CPU/PC[15] ), .I2(\CPU/PC[16] ), 
            .I3(\CPU/PC[17] ), .O(n1688)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2500.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2501 (.I0(n1658), .I1(n1659), .I2(n1660), .I3(n1688), 
            .O(n1689)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2501.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2502 (.I0(n1664), .I1(n1689), .I2(\CPU/PC[18] ), .O(n1690)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__2502.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__2503 (.I0(n1656), .I1(n623), .I2(n1665), .I3(\CPU/cycles[18] ), 
            .O(n1691)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2503.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2504 (.I0(\CPU/instr[18] ), .I1(n1666), .I2(n1690), 
            .I3(n1691), .O(n1692)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__2504.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__2505 (.I0(n1653), .I1(\mem_rdata[18] ), .I2(n1692), 
            .O(n1693)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2505.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2506 (.I0(n1640), .I1(n1687), .I2(n1693), .O(\CPU/writeBackData[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hefef */ ;
    defparam LUT__2506.LUTMASK = 16'hefef;
    EFX_LUT4 LUT__2507 (.I0(n1645), .I1(n1682), .I2(n683), .O(n1694)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__2507.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__2508 (.I0(n742), .I1(n681), .I2(n1694), .I3(n1646), 
            .O(n1695)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc355 */ ;
    defparam LUT__2508.LUTMASK = 16'hc355;
    EFX_LUT4 LUT__2509 (.I0(\CPU/rs2[19] ), .I1(\CPU/instr[31] ), .I2(\CPU/instr[4]~FF_frt_1_q ), 
            .I3(\CPU/instr[2]~FF_frt_0_q ), .O(n1549)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__2509.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__2510 (.I0(\CPU/instr[13] ), .I1(\CPU/instr[12] ), .I2(n1549), 
            .I3(\CPU/rs1[19] ), .O(n1696)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ccf */ ;
    defparam LUT__2510.LUTMASK = 16'h5ccf;
    EFX_LUT4 LUT__2511 (.I0(n1594), .I1(\CPU/aluReg[19] ), .I2(n1696), 
            .I3(\CPU/instr[14] ), .O(n1697)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077 */ ;
    defparam LUT__2511.LUTMASK = 16'h7077;
    EFX_LUT4 LUT__2512 (.I0(n1695), .I1(n1670), .I2(n1697), .I3(n1593), 
            .O(n1698)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__2512.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__2513 (.I0(n1689), .I1(\CPU/PC[18] ), .O(n1699)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2513.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2514 (.I0(n1664), .I1(n1699), .I2(\CPU/PC[19] ), .O(n1700)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__2514.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__2515 (.I0(\CPU/instr[19] ), .I1(n1666), .I2(n1665), 
            .I3(\CPU/cycles[19] ), .O(n1701)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2515.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2516 (.I0(n621), .I1(n1656), .I2(n1701), .O(n1702)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2516.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2517 (.I0(n1653), .I1(\mem_rdata[19] ), .I2(n1700), 
            .I3(n1702), .O(n1703)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__2517.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__2518 (.I0(n1640), .I1(n1698), .I2(n1703), .O(\CPU/writeBackData[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hefef */ ;
    defparam LUT__2518.LUTMASK = 16'hefef;
    EFX_LUT4 LUT__2519 (.I0(n1699), .I1(\CPU/PC[19] ), .I2(\CPU/PC[20] ), 
            .O(n1704)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__2519.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__2520 (.I0(n1608), .I1(n1621), .I2(\mult_dout[20] ), 
            .O(n1705)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__2520.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__2521 (.I0(n1609), .I1(\RAM_rdata[20] ), .I2(n1705), 
            .O(\mem_rdata[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__2521.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__2522 (.I0(n681), .I1(n683), .I2(n685), .I3(n687), 
            .O(n1706)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2522.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2523 (.I0(n1645), .I1(n1706), .I2(n679), .I3(n1646), 
            .O(n1707)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8700 */ ;
    defparam LUT__2523.LUTMASK = 16'h8700;
    EFX_LUT4 LUT__2524 (.I0(n1593), .I1(n1670), .O(n1708)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2524.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2525 (.I0(n740), .I1(n1646), .I2(n1708), .O(n1709)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__2525.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__2526 (.I0(\CPU/rs2[20] ), .I1(\CPU/instr[31] ), .I2(\CPU/instr[4]~FF_frt_1_q ), 
            .I3(\CPU/instr[2]~FF_frt_0_q ), .O(n1547)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__2526.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__2527 (.I0(\CPU/instr[13] ), .I1(\CPU/instr[12] ), .I2(n1547), 
            .I3(\CPU/rs1[20] ), .O(n1710)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ccf */ ;
    defparam LUT__2527.LUTMASK = 16'h5ccf;
    EFX_LUT4 LUT__2528 (.I0(n1593), .I1(\CPU/instr[14] ), .O(n1711)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2528.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2529 (.I0(n1710), .I1(n1711), .I2(n1707), .I3(n1709), 
            .O(n1712)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__2529.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__2530 (.I0(\CPU/instr[20] ), .I1(n1666), .I2(n1665), 
            .I3(\CPU/cycles[20] ), .O(n1713)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2530.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2531 (.I0(n1656), .I1(n619), .I2(n1595), .I3(\CPU/aluReg[20] ), 
            .O(n1714)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2531.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2532 (.I0(n1713), .I1(n1714), .O(n1715)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2532.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2533 (.I0(n1653), .I1(\mem_rdata[20] ), .I2(n1712), 
            .I3(n1715), .O(n1716)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7000 */ ;
    defparam LUT__2533.LUTMASK = 16'h7000;
    EFX_LUT4 LUT__2534 (.I0(n1664), .I1(n1704), .I2(n1640), .I3(n1716), 
            .O(\CPU/writeBackData[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4ff */ ;
    defparam LUT__2534.LUTMASK = 16'hf4ff;
    EFX_LUT4 LUT__2535 (.I0(n1645), .I1(n1706), .I2(n679), .I3(n677), 
            .O(n1717)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__2535.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__2536 (.I0(n738), .I1(n1717), .I2(n1646), .O(n1718)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__2536.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__2537 (.I0(\CPU/rs2[21] ), .I1(\CPU/instr[31] ), .I2(\CPU/instr[4]~FF_frt_1_q ), 
            .I3(\CPU/instr[2]~FF_frt_0_q ), .O(n1545)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__2537.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__2538 (.I0(\CPU/instr[13] ), .I1(\CPU/instr[12] ), .I2(n1545), 
            .I3(\CPU/rs1[21] ), .O(n1719)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ccf */ ;
    defparam LUT__2538.LUTMASK = 16'h5ccf;
    EFX_LUT4 LUT__2539 (.I0(n1594), .I1(\CPU/aluReg[21] ), .I2(n1719), 
            .I3(\CPU/instr[14] ), .O(n1720)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077 */ ;
    defparam LUT__2539.LUTMASK = 16'h7077;
    EFX_LUT4 LUT__2540 (.I0(n1718), .I1(n1670), .I2(n1720), .I3(n1593), 
            .O(n1721)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__2540.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__2541 (.I0(n1656), .I1(n617), .O(n1722)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2541.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2542 (.I0(n1622), .I1(\mult_dout[21] ), .I2(n1609), 
            .I3(\RAM_rdata[21] ), .O(\mem_rdata[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f88 */ ;
    defparam LUT__2542.LUTMASK = 16'h8f88;
    EFX_LUT4 LUT__2543 (.I0(\CPU/PC[19] ), .I1(\CPU/PC[20] ), .O(n1723)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2543.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2544 (.I0(n1699), .I1(n1723), .I2(n1664), .I3(\CPU/PC[21] ), 
            .O(n1724)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0708 */ ;
    defparam LUT__2544.LUTMASK = 16'h0708;
    EFX_LUT4 LUT__2545 (.I0(\CPU/instr[21] ), .I1(n1666), .I2(n1665), 
            .I3(\CPU/cycles[21] ), .O(n1725)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2545.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2546 (.I0(n1653), .I1(\mem_rdata[21] ), .I2(n1724), 
            .I3(n1725), .O(n1726)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__2546.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__2547 (.I0(n1640), .I1(n1721), .I2(n1722), .I3(n1726), 
            .O(\CPU/writeBackData[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfeff */ ;
    defparam LUT__2547.LUTMASK = 16'hfeff;
    EFX_LUT4 LUT__2548 (.I0(n1689), .I1(n1723), .I2(\CPU/PC[18] ), .I3(\CPU/PC[21] ), 
            .O(n1727)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2548.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2549 (.I0(n1727), .I1(\CPU/PC[22] ), .O(n1728)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__2549.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__2550 (.I0(n1664), .I1(n1728), .O(n1729)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2550.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2551 (.I0(n677), .I1(n679), .I2(n689), .I3(n691), 
            .O(n1730)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2551.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2552 (.I0(n1706), .I1(n1730), .O(n1731)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2552.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2553 (.I0(n6), .I1(n701), .O(n1732)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2553.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2554 (.I0(n1641), .I1(n1642), .I2(n1643), .I3(n1732), 
            .O(n1733)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2554.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2555 (.I0(n1731), .I1(n1733), .I2(n675), .O(n1734)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8787 */ ;
    defparam LUT__2555.LUTMASK = 16'h8787;
    EFX_LUT4 LUT__2556 (.I0(n736), .I1(n1734), .I2(n1646), .I3(n1708), 
            .O(n1735)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__2556.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__2557 (.I0(n1608), .I1(n1621), .I2(\mult_dout[22] ), 
            .O(n1736)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__2557.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__2558 (.I0(n1609), .I1(\RAM_rdata[22] ), .I2(n1736), 
            .O(\mem_rdata[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__2558.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__2559 (.I0(\CPU/rs2[22] ), .I1(\CPU/instr[31] ), .I2(\CPU/instr[4]~FF_frt_1_q ), 
            .I3(\CPU/instr[2]~FF_frt_0_q ), .O(n1543)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__2559.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__2560 (.I0(\CPU/instr[13] ), .I1(\CPU/instr[12] ), .I2(n1543), 
            .I3(\CPU/rs1[22] ), .O(n1737)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ccf */ ;
    defparam LUT__2560.LUTMASK = 16'h5ccf;
    EFX_LUT4 LUT__2561 (.I0(n1737), .I1(n1711), .O(n1738)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2561.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2562 (.I0(n1595), .I1(\CPU/aluReg[22] ), .O(n1739)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2562.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2563 (.I0(\CPU/instr[22] ), .I1(n1666), .I2(n1665), 
            .I3(\CPU/cycles[22] ), .O(n1740)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2563.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2564 (.I0(n615), .I1(n1656), .I2(n1739), .I3(n1740), 
            .O(n1741)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__2564.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__2565 (.I0(n1653), .I1(\mem_rdata[22] ), .I2(n1738), 
            .I3(n1741), .O(n1742)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__2565.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__2566 (.I0(n1640), .I1(n1729), .I2(n1735), .I3(n1742), 
            .O(\CPU/writeBackData[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfeff */ ;
    defparam LUT__2566.LUTMASK = 16'hfeff;
    EFX_LUT4 LUT__2567 (.I0(n1727), .I1(\CPU/PC[22] ), .I2(\CPU/PC[23] ), 
            .O(n1743)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__2567.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__2568 (.I0(n1731), .I1(n1733), .I2(n675), .O(n1744)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__2568.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__2569 (.I0(n734), .I1(n1646), .I2(n1708), .O(n1745)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__2569.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__2570 (.I0(n1646), .I1(n1744), .I2(n673), .I3(n1745), 
            .O(n1746)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7d00 */ ;
    defparam LUT__2570.LUTMASK = 16'h7d00;
    EFX_LUT4 LUT__2571 (.I0(n1609), .I1(\RAM_rdata[23] ), .I2(n1625), 
            .I3(n1653), .O(n1747)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__2571.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__2572 (.I0(\CPU/rs2[23] ), .I1(\CPU/instr[31] ), .I2(\CPU/instr[4]~FF_frt_1_q ), 
            .I3(\CPU/instr[2]~FF_frt_0_q ), .O(n1541)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__2572.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__2573 (.I0(\CPU/instr[13] ), .I1(\CPU/instr[12] ), .I2(n1541), 
            .I3(\CPU/rs1[23] ), .O(n1748)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ccf */ ;
    defparam LUT__2573.LUTMASK = 16'h5ccf;
    EFX_LUT4 LUT__2574 (.I0(n1748), .I1(n1711), .O(n1749)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2574.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2575 (.I0(n1595), .I1(\CPU/aluReg[23] ), .O(n1750)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2575.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2576 (.I0(n1656), .I1(n614), .I2(n1665), .I3(\CPU/cycles[23] ), 
            .O(n1751)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2576.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2577 (.I0(\CPU/instr[23] ), .I1(n1666), .I2(n1750), 
            .I3(n1751), .O(n1752)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__2577.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__2578 (.I0(n1746), .I1(n1747), .I2(n1749), .I3(n1752), 
            .O(n1753)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__2578.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__2579 (.I0(n1664), .I1(n1743), .I2(n1640), .I3(n1753), 
            .O(\CPU/writeBackData[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4ff */ ;
    defparam LUT__2579.LUTMASK = 16'hf4ff;
    EFX_LUT4 LUT__2580 (.I0(n1627), .I1(n1639), .I2(n1633), .O(n1754)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__2580.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__2581 (.I0(\CPU/instr[31] ), .I1(\CPU/rs2[24] ), .I2(\CPU/instr[4]~FF_frt_1_frt_2_q ), 
            .O(n1539)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__2581.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__2582 (.I0(\CPU/instr[13] ), .I1(\CPU/instr[12] ), .I2(n1539), 
            .I3(\CPU/rs1[24] ), .O(n1755)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ccf */ ;
    defparam LUT__2582.LUTMASK = 16'h5ccf;
    EFX_LUT4 LUT__2583 (.I0(n677), .I1(n679), .I2(n685), .I3(n687), 
            .O(n1756)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2583.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2584 (.I0(n673), .I1(n675), .O(n1757)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2584.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2585 (.I0(n1756), .I1(n1757), .I2(n681), .I3(n683), 
            .O(n1758)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2585.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2586 (.I0(n1645), .I1(n1758), .I2(n671), .I3(n1646), 
            .O(n1759)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8700 */ ;
    defparam LUT__2586.LUTMASK = 16'h8700;
    EFX_LUT4 LUT__2587 (.I0(n732), .I1(n1646), .I2(n1759), .I3(n1708), 
            .O(n1760)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__2587.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__2588 (.I0(\CPU/instr[24] ), .I1(n1666), .I2(n1665), 
            .I3(\CPU/cycles[24] ), .O(n1761)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2588.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2589 (.I0(\CPU/aluReg[24] ), .I1(n1595), .I2(n1761), 
            .O(n1762)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2589.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2590 (.I0(n1711), .I1(n1755), .I2(n1760), .I3(n1762), 
            .O(n1763)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__2590.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__2591 (.I0(n1622), .I1(\mult_dout[24] ), .I2(n1609), 
            .I3(\RAM_rdata[24] ), .O(\mem_rdata[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f88 */ ;
    defparam LUT__2591.LUTMASK = 16'h8f88;
    EFX_LUT4 LUT__2592 (.I0(n1754), .I1(n1763), .I2(\mem_rdata[24] ), 
            .I3(n1653), .O(\CPU/writeBackData[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0bb */ ;
    defparam LUT__2592.LUTMASK = 16'hf0bb;
    EFX_LUT4 LUT__2593 (.I0(\CPU/instr[31] ), .I1(\CPU/rs2[25] ), .I2(\CPU/instr[4]~FF_frt_1_frt_2_q ), 
            .O(n1537)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__2593.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__2594 (.I0(\CPU/instr[13] ), .I1(\CPU/instr[12] ), .I2(n1537), 
            .I3(\CPU/rs1[25] ), .O(n1764)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ccf */ ;
    defparam LUT__2594.LUTMASK = 16'h5ccf;
    EFX_LUT4 LUT__2595 (.I0(n673), .I1(n675), .I2(n677), .I3(n679), 
            .O(n1765)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2595.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2596 (.I0(n1706), .I1(n1765), .I2(n671), .I3(n1730), 
            .O(n1766)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2596.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2597 (.I0(n1733), .I1(n1766), .I2(n669), .I3(n1646), 
            .O(n1767)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8700 */ ;
    defparam LUT__2597.LUTMASK = 16'h8700;
    EFX_LUT4 LUT__2598 (.I0(n730), .I1(n1646), .I2(n1767), .I3(n1708), 
            .O(n1768)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__2598.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__2599 (.I0(\CPU/instr[25] ), .I1(n1666), .I2(n1665), 
            .I3(\CPU/cycles[25] ), .O(n1769)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2599.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2600 (.I0(\CPU/aluReg[25] ), .I1(n1595), .I2(n1769), 
            .O(n1770)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2600.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2601 (.I0(n1711), .I1(n1764), .I2(n1768), .I3(n1770), 
            .O(n1771)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__2601.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__2602 (.I0(n1622), .I1(\mult_dout[25] ), .I2(n1609), 
            .I3(\RAM_rdata[25] ), .O(\mem_rdata[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f88 */ ;
    defparam LUT__2602.LUTMASK = 16'h8f88;
    EFX_LUT4 LUT__2603 (.I0(n1754), .I1(n1771), .I2(\mem_rdata[25] ), 
            .I3(n1653), .O(\CPU/writeBackData[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0bb */ ;
    defparam LUT__2603.LUTMASK = 16'hf0bb;
    EFX_LUT4 LUT__2604 (.I0(n1622), .I1(\mult_dout[26] ), .I2(n1609), 
            .I3(\RAM_rdata[26] ), .O(\mem_rdata[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f88 */ ;
    defparam LUT__2604.LUTMASK = 16'h8f88;
    EFX_LUT4 LUT__2605 (.I0(\mem_rdata[26] ), .I1(n1653), .O(n1772)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2605.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2606 (.I0(n1733), .I1(n1766), .I2(n669), .O(n1773)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__2606.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__2607 (.I0(n728), .I1(n1646), .I2(n1708), .O(n1774)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__2607.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__2608 (.I0(n1646), .I1(n1773), .I2(n667), .I3(n1774), 
            .O(n1775)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7d00 */ ;
    defparam LUT__2608.LUTMASK = 16'h7d00;
    EFX_LUT4 LUT__2609 (.I0(\CPU/instr[31] ), .I1(\CPU/rs2[26] ), .I2(\CPU/instr[4]~FF_frt_1_frt_2_q ), 
            .O(n1535)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__2609.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__2610 (.I0(\CPU/instr[13] ), .I1(\CPU/instr[12] ), .I2(n1535), 
            .I3(\CPU/rs1[26] ), .O(n1776)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ccf */ ;
    defparam LUT__2610.LUTMASK = 16'h5ccf;
    EFX_LUT4 LUT__2611 (.I0(\CPU/cycles[26] ), .I1(n1665), .I2(n1595), 
            .I3(\CPU/aluReg[26] ), .O(n1777)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2611.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2612 (.I0(\CPU/instr[26] ), .I1(n1666), .I2(n1777), 
            .O(n1778)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2612.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2613 (.I0(n1711), .I1(n1776), .I2(n1778), .O(n1779)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__2613.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__2614 (.I0(n1640), .I1(n1772), .I2(n1775), .I3(n1779), 
            .O(\CPU/writeBackData[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfeff */ ;
    defparam LUT__2614.LUTMASK = 16'hfeff;
    EFX_LUT4 LUT__2616 (.I0(n1757), .I1(n667), .I2(n669), .I3(n671), 
            .O(n1781)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2616.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2367 (.I0(\mem_rdata[4] ), .I1(\mem_rdata[6] ), .O(n1588)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__2367.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__2617 (.I0(n1731), .I1(n1733), .I2(n1781), .O(n1782)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__2617.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__2618 (.I0(n1782), .I1(n665), .O(n1783)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__2618.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__2619 (.I0(n726), .I1(n1783), .I2(n1646), .I3(n1708), 
            .O(n1784)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__2619.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__2620 (.I0(\CPU/instr[31] ), .I1(\CPU/rs2[27] ), .I2(\CPU/instr[4]~FF_frt_1_frt_2_q ), 
            .O(n1533)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__2620.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__2621 (.I0(\CPU/instr[13] ), .I1(\CPU/instr[12] ), .I2(n1533), 
            .I3(\CPU/rs1[27] ), .O(n1785)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ccf */ ;
    defparam LUT__2621.LUTMASK = 16'h5ccf;
    EFX_LUT4 LUT__2622 (.I0(\CPU/cycles[27] ), .I1(n1665), .I2(n1595), 
            .I3(\CPU/aluReg[27] ), .O(n1786)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2622.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2623 (.I0(n1711), .I1(n1785), .I2(n1786), .O(n1787)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__2623.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__2624 (.I0(n1622), .I1(\mult_dout[27] ), .I2(n1609), 
            .I3(\RAM_rdata[27] ), .O(\mem_rdata[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f88 */ ;
    defparam LUT__2624.LUTMASK = 16'h8f88;
    EFX_LUT4 LUT__2625 (.I0(n1666), .I1(\CPU/instr[27] ), .I2(\mem_rdata[27] ), 
            .I3(n1653), .O(n1788)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2625.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2626 (.I0(n1640), .I1(n1784), .I2(n1787), .I3(n1788), 
            .O(\CPU/writeBackData[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hefff */ ;
    defparam LUT__2626.LUTMASK = 16'hefff;
    EFX_LUT4 LUT__2627 (.I0(n1782), .I1(n665), .I2(n663), .I3(n1646), 
            .O(n1789)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8700 */ ;
    defparam LUT__2627.LUTMASK = 16'h8700;
    EFX_LUT4 LUT__2628 (.I0(n724), .I1(n1646), .I2(n1789), .O(n1790)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__2628.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__2629 (.I0(n1622), .I1(\mult_dout[28] ), .I2(n1609), 
            .I3(\RAM_rdata[28] ), .O(\mem_rdata[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f88 */ ;
    defparam LUT__2629.LUTMASK = 16'h8f88;
    EFX_LUT4 LUT__2630 (.I0(\CPU/rs2[28] ), .I1(\CPU/instr[31] ), .I2(\CPU/instr[4]~FF_frt_1_q ), 
            .I3(\CPU/instr[2]~FF_frt_0_q ), .O(n1531)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__2630.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__2631 (.I0(\CPU/instr[13] ), .I1(\CPU/instr[12] ), .I2(n1531), 
            .I3(\CPU/rs1[28] ), .O(n1791)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ccf */ ;
    defparam LUT__2631.LUTMASK = 16'h5ccf;
    EFX_LUT4 LUT__2632 (.I0(n1791), .I1(n1711), .O(n1792)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2632.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2633 (.I0(\CPU/cycles[28] ), .I1(n1665), .I2(n1595), 
            .I3(\CPU/aluReg[28] ), .O(n1793)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2633.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2634 (.I0(\CPU/instr[28] ), .I1(n1666), .I2(n1793), 
            .O(n1794)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2634.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2635 (.I0(n1653), .I1(\mem_rdata[28] ), .I2(n1792), 
            .I3(n1794), .O(n1795)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__2635.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__2636 (.I0(n1708), .I1(n1790), .I2(n1640), .I3(n1795), 
            .O(\CPU/writeBackData[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8ff */ ;
    defparam LUT__2636.LUTMASK = 16'hf8ff;
    EFX_LUT4 LUT__2637 (.I0(n1782), .I1(n663), .I2(n665), .O(n1796)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__2637.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__2638 (.I0(n722), .I1(n661), .I2(n1796), .I3(n1646), 
            .O(n1797)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc355 */ ;
    defparam LUT__2638.LUTMASK = 16'hc355;
    EFX_LUT4 LUT__2639 (.I0(n1622), .I1(\mult_dout[29] ), .I2(n1609), 
            .I3(\RAM_rdata[29] ), .O(\mem_rdata[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f88 */ ;
    defparam LUT__2639.LUTMASK = 16'h8f88;
    EFX_LUT4 LUT__2640 (.I0(\CPU/rs2[29] ), .I1(\CPU/instr[31] ), .I2(\CPU/instr[4]~FF_frt_1_q ), 
            .I3(\CPU/instr[2]~FF_frt_0_q ), .O(n1529)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__2640.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__2641 (.I0(\CPU/instr[13] ), .I1(\CPU/instr[12] ), .I2(n1529), 
            .I3(\CPU/rs1[29] ), .O(n1798)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ccf */ ;
    defparam LUT__2641.LUTMASK = 16'h5ccf;
    EFX_LUT4 LUT__2642 (.I0(n1798), .I1(n1711), .O(n1799)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2642.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2643 (.I0(\CPU/instr[29] ), .I1(n1666), .I2(n1595), 
            .I3(\CPU/aluReg[29] ), .O(n1800)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2643.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2644 (.I0(\CPU/cycles[29] ), .I1(n1665), .I2(n1800), 
            .O(n1801)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2644.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2645 (.I0(n1653), .I1(\mem_rdata[29] ), .I2(n1799), 
            .I3(n1801), .O(n1802)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__2645.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__2646 (.I0(n1708), .I1(n1797), .I2(n1640), .I3(n1802), 
            .O(\CPU/writeBackData[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf2ff */ ;
    defparam LUT__2646.LUTMASK = 16'hf2ff;
    EFX_LUT4 LUT__2647 (.I0(n1796), .I1(n661), .I2(n659), .I3(n1646), 
            .O(n1803)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8700 */ ;
    defparam LUT__2647.LUTMASK = 16'h8700;
    EFX_LUT4 LUT__2648 (.I0(n720), .I1(n1646), .I2(n1708), .O(n1804)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__2648.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__2649 (.I0(n1622), .I1(\mult_dout[30] ), .I2(n1609), 
            .I3(\RAM_rdata[30] ), .O(\mem_rdata[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f88 */ ;
    defparam LUT__2649.LUTMASK = 16'h8f88;
    EFX_LUT4 LUT__2650 (.I0(\CPU/rs2[30] ), .I1(\CPU/instr[31] ), .I2(\CPU/instr[4]~FF_frt_1_q ), 
            .I3(\CPU/instr[2]~FF_frt_0_q ), .O(n1527)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__2650.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__2651 (.I0(\CPU/instr[13] ), .I1(\CPU/instr[12] ), .I2(n1527), 
            .I3(\CPU/rs1[30] ), .O(n1805)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ccf */ ;
    defparam LUT__2651.LUTMASK = 16'h5ccf;
    EFX_LUT4 LUT__2652 (.I0(n1805), .I1(n1711), .O(n1806)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2652.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2653 (.I0(\CPU/cycles[30] ), .I1(n1665), .I2(n1595), 
            .I3(\CPU/aluReg[30] ), .O(n1807)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2653.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2654 (.I0(\CPU/instr[30] ), .I1(n1666), .I2(n1807), 
            .O(n1808)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2654.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2655 (.I0(n1653), .I1(\mem_rdata[30] ), .I2(n1806), 
            .I3(n1808), .O(n1809)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__2655.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__2656 (.I0(n1804), .I1(n1803), .I2(n1640), .I3(n1809), 
            .O(\CPU/writeBackData[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf2ff */ ;
    defparam LUT__2656.LUTMASK = 16'hf2ff;
    EFX_LUT4 LUT__2657 (.I0(n659), .I1(n661), .I2(n663), .I3(n665), 
            .O(n1810)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2657.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2658 (.I0(n1731), .I1(n1733), .I2(n1781), .I3(n1810), 
            .O(n1811)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2658.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2659 (.I0(n719), .I1(n657), .I2(n1811), .I3(n1646), 
            .O(n1812)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc355 */ ;
    defparam LUT__2659.LUTMASK = 16'hc355;
    EFX_LUT4 LUT__2660 (.I0(\CPU/rs2[31] ), .I1(\CPU/instr[31] ), .I2(\CPU/instr[4]~FF_frt_1_q ), 
            .I3(\CPU/instr[2]~FF_frt_0_q ), .O(n1525)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__2660.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__2661 (.I0(n1649), .I1(n1673), .I2(n1525), .I3(\CPU/rs1[31] ), 
            .O(n1813)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h533f */ ;
    defparam LUT__2661.LUTMASK = 16'h533f;
    EFX_LUT4 LUT__2662 (.I0(\CPU/aluReg[31] ), .I1(n1594), .I2(n1813), 
            .O(n1814)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2662.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2663 (.I0(n1812), .I1(n1670), .I2(n1814), .I3(n1593), 
            .O(n1815)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__2663.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__2664 (.I0(n1622), .I1(\mult_dout[31] ), .I2(n1630), 
            .O(\mem_rdata[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8 */ ;
    defparam LUT__2664.LUTMASK = 16'hf8f8;
    EFX_LUT4 LUT__2665 (.I0(\CPU/instr[31] ), .I1(n1666), .I2(n1665), 
            .I3(\CPU/cycles[31] ), .O(n1816)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2665.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2666 (.I0(n1653), .I1(\mem_rdata[31] ), .I2(n1816), 
            .O(n1817)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__2666.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__2667 (.I0(n1640), .I1(n1815), .I2(n1817), .O(\CPU/writeBackData[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hefef */ ;
    defparam LUT__2667.LUTMASK = 16'hefef;
    EFX_LUT4 LUT__2668 (.I0(\CPU/instr[7] ), .I1(\CPU/instr[8] ), .I2(\CPU/instr[9] ), 
            .I3(\CPU/instr[10] ), .O(n1818)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__2668.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__2669 (.I0(\CPU/instr[11] ), .I1(n1818), .O(\CPU/not_equal_22/n9 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__2669.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__2670 (.I0(\CPU/state[3] ), .I1(\CPU/state[2] ), .I2(\CPU/instr[4] ), 
            .I3(\CPU/instr[2]~FF_frt_0_q ), .O(\CPU/writeBack )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0ee */ ;
    defparam LUT__2670.LUTMASK = 16'he0ee;
    EFX_LUT4 LUT__2671 (.I0(n1608), .I1(n1621), .I2(\mult_dout[8] ), .O(n1819)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__2671.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__2672 (.I0(n1603), .I1(n1602), .I2(n1608), .I3(\RAM_rdata[8] ), 
            .O(n1820)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__2672.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__2673 (.I0(n1600), .I1(n1614), .I2(n1608), .I3(\uart_dout[8] ), 
            .O(n1821)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__2673.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__2674 (.I0(n1819), .I1(n1820), .I2(n1821), .O(\mem_rdata[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfefe */ ;
    defparam LUT__2674.LUTMASK = 16'hfefe;
    EFX_LUT4 LUT__2675 (.I0(\CPU/instr[12] ), .I1(n12), .O(n1822)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2675.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2676 (.I0(\CPU/instr[13] ), .I1(n1822), .O(n1823)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2676.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2677 (.I0(\mem_rdata[8] ), .I1(\mem_rdata[24] ), .I2(n612), 
            .I3(n1823), .O(n1824)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__2677.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__2678 (.I0(\CPU/instr[13] ), .I1(n612), .O(n1825)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2678.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2679 (.I0(n1822), .I1(n1825), .O(n1826)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2679.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2680 (.I0(n1608), .I1(n1621), .I2(\mult_dout[0] ), .O(n1827)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__2680.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__2681 (.I0(n1600), .I1(n1614), .I2(n1608), .I3(\uart_dout[0] ), 
            .O(n1828)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__2681.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__2682 (.I0(n1603), .I1(n1602), .I2(n1608), .I3(\RAM_rdata[0] ), 
            .O(n1829)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__2682.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__2683 (.I0(n1823), .I1(n1825), .O(n1830)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__2683.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__2684 (.I0(n1827), .I1(n1828), .I2(n1829), .I3(n1830), 
            .O(n1831)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__2684.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__2685 (.I0(n1826), .I1(\mem_rdata[16] ), .I2(n1831), 
            .I3(n1599), .O(n1832)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__2685.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__2686 (.I0(\CPU/rs1[31] ), .I1(\CPU/instr[12] ), .I2(n1525), 
            .O(n1833)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__2686.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__2687 (.I0(n657), .I1(n667), .I2(n669), .I3(n671), 
            .O(n1834)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2687.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2688 (.I0(n1706), .I1(n1765), .I2(n1810), .I3(n1834), 
            .O(n1835)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2688.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2689 (.I0(n1645), .I1(n1835), .I2(n658), .O(n1836)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__2689.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__2690 (.I0(n1525), .I1(\CPU/instr[12] ), .I2(\CPU/rs1[31] ), 
            .I3(\CPU/instr[14] ), .O(n1837)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__2690.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__2691 (.I0(\CPU/rs1[0] ), .I1(n1587), .I2(\CPU/instr[14] ), 
            .I3(\CPU/instr[13] ), .O(n1838)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__2691.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__2692 (.I0(n1836), .I1(n1833), .I2(n1837), .I3(n1838), 
            .O(n1839)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__2692.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__2693 (.I0(n1587), .I1(\CPU/rs1[0] ), .I2(n1673), .O(n1840)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__2693.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__2694 (.I0(n780), .I1(n6), .I2(n1646), .I3(n1670), 
            .O(n1841)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__2694.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__2695 (.I0(\CPU/aluReg[0] ), .I1(n1594), .I2(n1840), 
            .I3(n1841), .O(n1842)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__2695.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__2696 (.I0(n1842), .I1(n1839), .I2(n1593), .O(n1843)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__2696.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__2697 (.I0(n1665), .I1(\CPU/cycles[0] ), .O(n1844)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2697.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2698 (.I0(n1832), .I1(n1824), .I2(n1843), .I3(n1844), 
            .O(\CPU/writeBackData[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff2 */ ;
    defparam LUT__2698.LUTMASK = 16'hfff2;
    EFX_LUT4 LUT__2699 (.I0(n1603), .I1(n1602), .I2(n1608), .I3(\RAM_rdata[9] ), 
            .O(n1845)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__2699.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__2700 (.I0(n1608), .I1(n1621), .I2(\mult_dout[9] ), .O(n1846)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__2700.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__2701 (.I0(n1600), .I1(n1614), .I2(n1608), .I3(\uart_dout[9] ), 
            .O(n1847)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__2701.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__2702 (.I0(n1845), .I1(n1846), .I2(n1847), .O(\mem_rdata[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfefe */ ;
    defparam LUT__2702.LUTMASK = 16'hfefe;
    EFX_LUT4 LUT__2703 (.I0(\mem_rdata[9] ), .I1(\mem_rdata[25] ), .I2(n612), 
            .I3(n1823), .O(n1848)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__2703.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__2704 (.I0(n1608), .I1(n1621), .I2(\mult_dout[1] ), .O(n1849)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__2704.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__2705 (.I0(n1600), .I1(n1614), .I2(n1608), .I3(\uart_dout[1] ), 
            .O(n1850)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__2705.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__2706 (.I0(n1603), .I1(n1602), .I2(n1608), .I3(\RAM_rdata[1] ), 
            .O(n1851)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__2706.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__2707 (.I0(n1849), .I1(n1850), .I2(n1851), .I3(n1830), 
            .O(n1852)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__2707.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__2708 (.I0(n1826), .I1(\mem_rdata[17] ), .I2(n1852), 
            .I3(n1599), .O(n1853)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__2708.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__2709 (.I0(\mem_wdata[1] ), .I1(\CPU/instr[21] ), .I2(\CPU/instr[4]~FF_frt_1_q ), 
            .I3(\CPU/instr[2]~FF_frt_0_q ), .O(n1585)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__2709.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__2710 (.I0(\CPU/instr[13] ), .I1(\CPU/instr[12] ), .I2(n1585), 
            .I3(\CPU/rs1[1] ), .O(n1854)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ccf */ ;
    defparam LUT__2710.LUTMASK = 16'h5ccf;
    EFX_LUT4 LUT__2711 (.I0(n778), .I1(n6), .I2(n717), .I3(n1646), .O(n1855)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc355 */ ;
    defparam LUT__2711.LUTMASK = 16'hc355;
    EFX_LUT4 LUT__2712 (.I0(n1594), .I1(\CPU/aluReg[1] ), .I2(n1855), 
            .I3(n1670), .O(n1856)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077 */ ;
    defparam LUT__2712.LUTMASK = 16'h7077;
    EFX_LUT4 LUT__2713 (.I0(n1854), .I1(\CPU/instr[14] ), .I2(n1856), 
            .I3(n1593), .O(n1857)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__2713.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__2714 (.I0(n8), .I1(n1656), .I2(n1664), .I3(\CPU/PC[1] ), 
            .O(n1858)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077 */ ;
    defparam LUT__2714.LUTMASK = 16'h7077;
    EFX_LUT4 LUT__2715 (.I0(\CPU/cycles[1] ), .I1(n1665), .I2(n1857), 
            .I3(n1858), .O(n1859)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__2715.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__2716 (.I0(n1848), .I1(n1853), .I2(n1859), .O(\CPU/writeBackData[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f */ ;
    defparam LUT__2716.LUTMASK = 16'h4f4f;
    EFX_LUT4 LUT__2717 (.I0(n1622), .I1(\mult_dout[10] ), .I2(n1609), 
            .I3(\RAM_rdata[10] ), .O(\mem_rdata[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f88 */ ;
    defparam LUT__2717.LUTMASK = 16'h8f88;
    EFX_LUT4 LUT__2718 (.I0(\mem_rdata[10] ), .I1(\mem_rdata[26] ), .I2(n612), 
            .I3(n1823), .O(n1860)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__2718.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__2719 (.I0(n1600), .I1(n1614), .I2(n1608), .O(n1861)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__2719.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__2720 (.I0(n1603), .I1(n1602), .I2(n1608), .I3(\RAM_rdata[2] ), 
            .O(n1862)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__2720.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__2721 (.I0(n1608), .I1(n1621), .I2(\mult_dout[2] ), .O(n1863)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__2721.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__2722 (.I0(\uart_dout[2] ), .I1(n1861), .I2(n1862), .I3(n1863), 
            .O(\mem_rdata[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8 */ ;
    defparam LUT__2722.LUTMASK = 16'hfff8;
    EFX_LUT4 LUT__2723 (.I0(\mem_rdata[2] ), .I1(n1830), .I2(\mem_rdata[18] ), 
            .I3(n1826), .O(n1864)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__2723.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__2724 (.I0(\mem_wdata[2] ), .I1(\CPU/instr[22] ), .I2(\CPU/instr[4]~FF_frt_1_q ), 
            .I3(\CPU/instr[2]~FF_frt_0_q ), .O(n1583)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__2724.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__2725 (.I0(\CPU/instr[13] ), .I1(\CPU/instr[12] ), .I2(n1583), 
            .I3(\CPU/rs1[2] ), .O(n1865)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ccf */ ;
    defparam LUT__2725.LUTMASK = 16'h5ccf;
    EFX_LUT4 LUT__2726 (.I0(n6), .I1(n717), .O(n1866)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2726.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2727 (.I0(n776), .I1(n1866), .I2(n715), .I3(n1646), 
            .O(n1867)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc355 */ ;
    defparam LUT__2727.LUTMASK = 16'hc355;
    EFX_LUT4 LUT__2728 (.I0(n1594), .I1(\CPU/aluReg[2] ), .I2(n1867), 
            .I3(n1670), .O(n1868)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077 */ ;
    defparam LUT__2728.LUTMASK = 16'h7077;
    EFX_LUT4 LUT__2729 (.I0(n1865), .I1(\CPU/instr[14] ), .I2(n1868), 
            .I3(n1593), .O(n1869)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__2729.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__2730 (.I0(n1656), .I1(n655), .I2(n1665), .I3(\CPU/cycles[2] ), 
            .O(n1870)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2730.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2731 (.I0(\CPU/PC[2] ), .I1(n1664), .I2(n1869), .I3(n1870), 
            .O(n1871)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__2731.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__2732 (.I0(n1860), .I1(n1864), .I2(n1599), .I3(n1871), 
            .O(\CPU/writeBackData[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h40ff */ ;
    defparam LUT__2732.LUTMASK = 16'h40ff;
    EFX_LUT4 LUT__2733 (.I0(n1622), .I1(\mult_dout[11] ), .I2(n1609), 
            .I3(\RAM_rdata[11] ), .O(\mem_rdata[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f88 */ ;
    defparam LUT__2733.LUTMASK = 16'h8f88;
    EFX_LUT4 LUT__2734 (.I0(\mem_rdata[11] ), .I1(\mem_rdata[27] ), .I2(n612), 
            .I3(n1823), .O(n1872)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__2734.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__2735 (.I0(n1603), .I1(n1602), .I2(n1608), .I3(\RAM_rdata[3] ), 
            .O(n1873)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__2735.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__2736 (.I0(n1608), .I1(n1621), .I2(\mult_dout[3] ), .O(n1874)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__2736.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__2737 (.I0(\uart_dout[3] ), .I1(n1861), .I2(n1873), .I3(n1874), 
            .O(\mem_rdata[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8 */ ;
    defparam LUT__2737.LUTMASK = 16'hfff8;
    EFX_LUT4 LUT__2738 (.I0(\RAM_rdata[19] ), .I1(n1609), .I2(n1624), 
            .I3(n1826), .O(n1875)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__2738.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__2739 (.I0(n1830), .I1(\mem_rdata[3] ), .I2(n1875), .I3(n1599), 
            .O(n1876)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__2739.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__2740 (.I0(n1866), .I1(n715), .I2(n713), .O(n1877)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__2740.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__2741 (.I0(n774), .I1(n1877), .I2(\CPU/instr[13] ), .I3(n1646), 
            .O(n1878)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__2741.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__2742 (.I0(\mem_wdata[3] ), .I1(\CPU/instr[23] ), .I2(\CPU/instr[4]~FF_frt_1_frt_2_q ), 
            .I3(\CPU/rs1[3] ), .O(n1879)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac53 */ ;
    defparam LUT__2742.LUTMASK = 16'hac53;
    EFX_LUT4 LUT__2743 (.I0(n1879), .I1(n1878), .I2(\CPU/instr[12] ), 
            .I3(\CPU/instr[14] ), .O(n1880)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h050c */ ;
    defparam LUT__2743.LUTMASK = 16'h050c;
    EFX_LUT4 LUT__2744 (.I0(\CPU/instr[23] ), .I1(\mem_wdata[3] ), .I2(\CPU/instr[4]~FF_frt_1_frt_2_q ), 
            .O(n1581)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__2744.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__2745 (.I0(n1594), .I1(\CPU/aluReg[3] ), .O(n1881)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2745.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2746 (.I0(\CPU/rs1[3] ), .I1(n1649), .I2(n1581), .I3(n1881), 
            .O(n1882)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007f */ ;
    defparam LUT__2746.LUTMASK = 16'h007f;
    EFX_LUT4 LUT__2747 (.I0(n1882), .I1(n1880), .I2(n1593), .O(n1883)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__2747.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__2748 (.I0(\CPU/PC[2] ), .I1(\CPU/PC[3] ), .O(n1884)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__2748.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__2749 (.I0(n1656), .I1(n653), .I2(n1665), .I3(\CPU/cycles[3] ), 
            .O(n1885)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2749.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2750 (.I0(n1884), .I1(n1664), .I2(n1885), .O(n1886)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__2750.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__2751 (.I0(n1876), .I1(n1872), .I2(n1883), .I3(n1886), 
            .O(\CPU/writeBackData[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf2ff */ ;
    defparam LUT__2751.LUTMASK = 16'hf2ff;
    EFX_LUT4 LUT__2752 (.I0(n1622), .I1(\mult_dout[12] ), .I2(n1609), 
            .I3(\RAM_rdata[12] ), .O(\mem_rdata[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f88 */ ;
    defparam LUT__2752.LUTMASK = 16'h8f88;
    EFX_LUT4 LUT__2753 (.I0(\mem_rdata[12] ), .I1(\mem_rdata[28] ), .I2(n612), 
            .I3(n1823), .O(n1887)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__2753.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__2754 (.I0(n1600), .I1(n1614), .I2(n1608), .I3(\uart_dout[4] ), 
            .O(n1888)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__2754.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__2755 (.I0(n1608), .I1(n1621), .I2(\mult_dout[4] ), .O(n1889)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__2755.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__2756 (.I0(\RAM_rdata[4] ), .I1(n1609), .I2(n1888), .I3(n1889), 
            .O(\mem_rdata[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff2 */ ;
    defparam LUT__2756.LUTMASK = 16'hfff2;
    EFX_LUT4 LUT__2757 (.I0(\mem_rdata[4] ), .I1(n1830), .I2(\mem_rdata[20] ), 
            .I3(n1826), .O(n1890)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__2757.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__2758 (.I0(\CPU/PC[2] ), .I1(\CPU/PC[3] ), .I2(\CPU/PC[4] ), 
            .O(n1891)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8787 */ ;
    defparam LUT__2758.LUTMASK = 16'h8787;
    EFX_LUT4 LUT__2759 (.I0(\mem_wdata[4] ), .I1(\CPU/instr[24] ), .I2(\CPU/instr[4]~FF_frt_1_q ), 
            .I3(\CPU/instr[2]~FF_frt_0_q ), .O(n1579)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__2759.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__2760 (.I0(\CPU/instr[13] ), .I1(\CPU/instr[12] ), .I2(n1579), 
            .I3(\CPU/rs1[4] ), .O(n1892)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ccf */ ;
    defparam LUT__2760.LUTMASK = 16'h5ccf;
    EFX_LUT4 LUT__2761 (.I0(n6), .I1(n713), .I2(n715), .I3(n717), .O(n1893)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2761.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2762 (.I0(n772), .I1(n1893), .I2(n711), .I3(n1646), 
            .O(n1894)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc355 */ ;
    defparam LUT__2762.LUTMASK = 16'hc355;
    EFX_LUT4 LUT__2763 (.I0(n1594), .I1(\CPU/aluReg[4] ), .I2(n1894), 
            .I3(n1670), .O(n1895)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077 */ ;
    defparam LUT__2763.LUTMASK = 16'h7077;
    EFX_LUT4 LUT__2764 (.I0(n1892), .I1(\CPU/instr[14] ), .I2(n1895), 
            .I3(n1593), .O(n1896)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__2764.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__2765 (.I0(n1656), .I1(n651), .I2(n1665), .I3(\CPU/cycles[4] ), 
            .O(n1897)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2765.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2766 (.I0(n1891), .I1(n1664), .I2(n1896), .I3(n1897), 
            .O(n1898)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__2766.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__2767 (.I0(n1887), .I1(n1890), .I2(n1599), .I3(n1898), 
            .O(\CPU/writeBackData[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h40ff */ ;
    defparam LUT__2767.LUTMASK = 16'h40ff;
    EFX_LUT4 LUT__2768 (.I0(n1622), .I1(\mult_dout[13] ), .I2(n1609), 
            .I3(\RAM_rdata[13] ), .O(\mem_rdata[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f88 */ ;
    defparam LUT__2768.LUTMASK = 16'h8f88;
    EFX_LUT4 LUT__2769 (.I0(\mem_rdata[13] ), .I1(\mem_rdata[29] ), .I2(n612), 
            .I3(n1823), .O(n1899)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__2769.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__2770 (.I0(n1600), .I1(n1614), .I2(n1608), .I3(\uart_dout[5] ), 
            .O(n1900)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__2770.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__2771 (.I0(n1608), .I1(n1621), .I2(\mult_dout[5] ), .O(n1901)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__2771.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__2772 (.I0(\RAM_rdata[5] ), .I1(n1609), .I2(n1900), .I3(n1901), 
            .O(\mem_rdata[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff2 */ ;
    defparam LUT__2772.LUTMASK = 16'hfff2;
    EFX_LUT4 LUT__2773 (.I0(\mem_rdata[5] ), .I1(n1830), .I2(\mem_rdata[21] ), 
            .I3(n1826), .O(n1902)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__2773.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__2774 (.I0(\CPU/PC[2] ), .I1(\CPU/PC[3] ), .I2(\CPU/PC[4] ), 
            .I3(\CPU/PC[5] ), .O(n1903)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h807f */ ;
    defparam LUT__2774.LUTMASK = 16'h807f;
    EFX_LUT4 LUT__2775 (.I0(\mem_wdata[5] ), .I1(\CPU/instr[25] ), .I2(\CPU/instr[4]~FF_frt_1_q ), 
            .I3(\CPU/instr[2]~FF_frt_0_q ), .O(n1577)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__2775.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__2776 (.I0(\CPU/instr[13] ), .I1(\CPU/instr[12] ), .I2(n1577), 
            .I3(\CPU/rs1[5] ), .O(n1904)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ccf */ ;
    defparam LUT__2776.LUTMASK = 16'h5ccf;
    EFX_LUT4 LUT__2777 (.I0(n1893), .I1(n711), .I2(n709), .I3(n1646), 
            .O(n1905)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8700 */ ;
    defparam LUT__2777.LUTMASK = 16'h8700;
    EFX_LUT4 LUT__2778 (.I0(n770), .I1(n1646), .I2(n1670), .O(n1906)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__2778.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__2779 (.I0(n1594), .I1(\CPU/aluReg[5] ), .I2(n1905), 
            .I3(n1906), .O(n1907)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077 */ ;
    defparam LUT__2779.LUTMASK = 16'h7077;
    EFX_LUT4 LUT__2780 (.I0(n1904), .I1(\CPU/instr[14] ), .I2(n1907), 
            .I3(n1593), .O(n1908)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__2780.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__2781 (.I0(n1656), .I1(n649), .I2(n1665), .I3(\CPU/cycles[5] ), 
            .O(n1909)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2781.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2782 (.I0(n1903), .I1(n1664), .I2(n1908), .I3(n1909), 
            .O(n1910)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__2782.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__2783 (.I0(n1899), .I1(n1902), .I2(n1599), .I3(n1910), 
            .O(\CPU/writeBackData[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h40ff */ ;
    defparam LUT__2783.LUTMASK = 16'h40ff;
    EFX_LUT4 LUT__2784 (.I0(n1622), .I1(\mult_dout[14] ), .I2(n1609), 
            .I3(\RAM_rdata[14] ), .O(\mem_rdata[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f88 */ ;
    defparam LUT__2784.LUTMASK = 16'h8f88;
    EFX_LUT4 LUT__2785 (.I0(\mem_rdata[14] ), .I1(\mem_rdata[30] ), .I2(n612), 
            .I3(n1823), .O(n1911)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__2785.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__2786 (.I0(n1603), .I1(n1602), .I2(n1608), .I3(\RAM_rdata[6] ), 
            .O(n1912)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__2786.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__2787 (.I0(n1608), .I1(n1621), .I2(\mult_dout[6] ), .O(n1913)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__2787.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__2788 (.I0(\uart_dout[6] ), .I1(n1861), .I2(n1912), .I3(n1913), 
            .O(\mem_rdata[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8 */ ;
    defparam LUT__2788.LUTMASK = 16'hfff8;
    EFX_LUT4 LUT__2789 (.I0(\RAM_rdata[22] ), .I1(n1609), .I2(n1736), 
            .I3(n1826), .O(n1914)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__2789.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__2790 (.I0(n1830), .I1(\mem_rdata[6] ), .I2(n1914), .I3(n1599), 
            .O(n1915)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__2790.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__2791 (.I0(n1656), .I1(n647), .O(n1916)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2791.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2792 (.I0(\mem_wdata[6] ), .I1(\CPU/instr[26] ), .I2(\CPU/instr[4]~FF_frt_1_q ), 
            .I3(\CPU/instr[2]~FF_frt_0_q ), .O(n1575)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__2792.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__2793 (.I0(n1649), .I1(n1673), .I2(\CPU/rs1[6] ), .I3(n1575), 
            .O(n1917)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h533f */ ;
    defparam LUT__2793.LUTMASK = 16'h533f;
    EFX_LUT4 LUT__2794 (.I0(n1642), .I1(n1866), .I2(n707), .I3(n1646), 
            .O(n1918)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8700 */ ;
    defparam LUT__2794.LUTMASK = 16'h8700;
    EFX_LUT4 LUT__2795 (.I0(n768), .I1(n1646), .I2(n1918), .I3(n1670), 
            .O(n1919)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__2795.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__2796 (.I0(n1594), .I1(\CPU/aluReg[6] ), .O(n1920)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2796.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2797 (.I0(n1919), .I1(n1920), .I2(n1917), .I3(n1593), 
            .O(n1921)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__2797.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__2798 (.I0(n1658), .I1(\CPU/PC[6] ), .O(n1922)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__2798.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__2799 (.I0(n1664), .I1(n1922), .O(n1923)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__2799.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__2800 (.I0(\CPU/cycles[6] ), .I1(n1665), .I2(n1921), 
            .I3(n1923), .O(n1924)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__2800.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__2801 (.I0(n1915), .I1(n1911), .I2(n1916), .I3(n1924), 
            .O(\CPU/writeBackData[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf2ff */ ;
    defparam LUT__2801.LUTMASK = 16'hf2ff;
    EFX_LUT4 LUT__2802 (.I0(\mem_rdata[31] ), .I1(\mem_rdata[15] ), .I2(n612), 
            .I3(n1822), .O(n1925)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__2802.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__2803 (.I0(n1609), .I1(\RAM_rdata[23] ), .I2(n1625), 
            .O(\mem_rdata[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__2803.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__2804 (.I0(n1634), .I1(n1636), .O(\mem_rdata[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__2804.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__2805 (.I0(\mem_rdata[7] ), .I1(\mem_rdata[23] ), .I2(n1822), 
            .I3(n612), .O(n1926)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__2805.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__2806 (.I0(\CPU/instr[13] ), .I1(n1599), .O(n1927)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2806.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2807 (.I0(\mem_wdata[7] ), .I1(\CPU/instr[27] ), .I2(\CPU/instr[4]~FF_frt_1_q ), 
            .I3(\CPU/instr[2]~FF_frt_0_q ), .O(n1573)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__2807.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__2808 (.I0(\CPU/instr[13] ), .I1(\CPU/instr[12] ), .I2(n1573), 
            .I3(\CPU/rs1[7] ), .O(n1928)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ccf */ ;
    defparam LUT__2808.LUTMASK = 16'h5ccf;
    EFX_LUT4 LUT__2809 (.I0(n6), .I1(n707), .I2(n717), .O(n1929)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__2809.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__2810 (.I0(n1642), .I1(n1929), .I2(n705), .I3(n1646), 
            .O(n1930)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8700 */ ;
    defparam LUT__2810.LUTMASK = 16'h8700;
    EFX_LUT4 LUT__2811 (.I0(n766), .I1(n1646), .I2(n1670), .O(n1931)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__2811.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__2812 (.I0(n1594), .I1(\CPU/aluReg[7] ), .I2(n1930), 
            .I3(n1931), .O(n1932)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077 */ ;
    defparam LUT__2812.LUTMASK = 16'h7077;
    EFX_LUT4 LUT__2813 (.I0(n1928), .I1(\CPU/instr[14] ), .I2(n1932), 
            .I3(n1593), .O(n1933)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__2813.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__2814 (.I0(n1658), .I1(\CPU/PC[6] ), .I2(\CPU/PC[7] ), 
            .O(n1934)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8787 */ ;
    defparam LUT__2814.LUTMASK = 16'h8787;
    EFX_LUT4 LUT__2815 (.I0(n1656), .I1(n645), .I2(n1665), .I3(\CPU/cycles[7] ), 
            .O(n1935)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2815.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2816 (.I0(n1934), .I1(n1664), .I2(n1935), .O(n1936)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__2816.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__2817 (.I0(n1653), .I1(\mem_rdata[7] ), .I2(n1933), .I3(n1936), 
            .O(n1937)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__2817.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__2818 (.I0(n1926), .I1(n1925), .I2(n1927), .I3(n1937), 
            .O(\CPU/writeBackData[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0ff */ ;
    defparam LUT__2818.LUTMASK = 16'he0ff;
    EFX_LUT4 LUT__2819 (.I0(\mem_rdata[8] ), .I1(\CPU/instr[13] ), .O(n1938)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2819.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2820 (.I0(n1611), .I1(n1599), .O(n1939)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2820.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2821 (.I0(n1627), .I1(n1633), .I2(n1639), .I3(n1939), 
            .O(n1940)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf */ ;
    defparam LUT__2821.LUTMASK = 16'h00bf;
    EFX_LUT4 LUT__2822 (.I0(\mem_rdata[24] ), .I1(\mem_rdata[8] ), .I2(n1825), 
            .I3(\CPU/instr[12] ), .O(n1941)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__2822.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__2823 (.I0(\CPU/rs2[8] ), .I1(\CPU/instr[28] ), .I2(\CPU/instr[4]~FF_frt_1_q ), 
            .I3(\CPU/instr[2]~FF_frt_0_q ), .O(n1571)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__2823.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__2824 (.I0(\CPU/instr[13] ), .I1(\CPU/instr[12] ), .I2(n1571), 
            .I3(\CPU/rs1[8] ), .O(n1942)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ccf */ ;
    defparam LUT__2824.LUTMASK = 16'h5ccf;
    EFX_LUT4 LUT__2825 (.I0(n1594), .I1(\CPU/aluReg[8] ), .O(n1943)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2825.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2826 (.I0(n6), .I1(n705), .I2(n707), .I3(n717), .O(n1944)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2826.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2827 (.I0(n1642), .I1(n1944), .I2(n703), .I3(n1646), 
            .O(n1945)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8700 */ ;
    defparam LUT__2827.LUTMASK = 16'h8700;
    EFX_LUT4 LUT__2828 (.I0(n764), .I1(n1646), .I2(n1945), .I3(n1670), 
            .O(n1946)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__2828.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__2829 (.I0(\CPU/instr[14] ), .I1(n1942), .I2(n1943), 
            .I3(n1946), .O(n1947)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__2829.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__2830 (.I0(\CPU/PC[6] ), .I1(\CPU/PC[7] ), .O(n1948)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2830.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2831 (.I0(n1658), .I1(n1948), .O(n1949)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2831.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2832 (.I0(n1949), .I1(\CPU/PC[8] ), .O(n1950)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__2832.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__2833 (.I0(n1656), .I1(n643), .I2(n1665), .I3(\CPU/cycles[8] ), 
            .O(n1951)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2833.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2834 (.I0(n1664), .I1(n1950), .I2(n1951), .O(n1952)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__2834.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__2835 (.I0(n1593), .I1(n1947), .I2(n1952), .O(n1953)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__2835.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__2836 (.I0(n1940), .I1(n1941), .I2(n1938), .I3(n1953), 
            .O(\CPU/writeBackData[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h01ff */ ;
    defparam LUT__2836.LUTMASK = 16'h01ff;
    EFX_LUT4 LUT__2837 (.I0(\mem_rdata[9] ), .I1(\CPU/instr[13] ), .O(n1954)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2837.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2838 (.I0(\mem_rdata[25] ), .I1(\mem_rdata[9] ), .I2(n1825), 
            .I3(\CPU/instr[12] ), .O(n1955)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__2838.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__2839 (.I0(n1949), .I1(\CPU/PC[8] ), .I2(\CPU/PC[9] ), 
            .O(n1956)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8787 */ ;
    defparam LUT__2839.LUTMASK = 16'h8787;
    EFX_LUT4 LUT__2840 (.I0(n1664), .I1(n1956), .O(n1957)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__2840.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__2841 (.I0(n1595), .I1(\CPU/aluReg[9] ), .O(n1958)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2841.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2842 (.I0(\CPU/rs2[9] ), .I1(\CPU/instr[29] ), .I2(\CPU/instr[4]~FF_frt_1_q ), 
            .I3(\CPU/instr[2]~FF_frt_0_q ), .O(n1569)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__2842.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__2843 (.I0(\CPU/instr[13] ), .I1(\CPU/instr[12] ), .I2(n1569), 
            .I3(\CPU/rs1[9] ), .O(n1959)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ccf */ ;
    defparam LUT__2843.LUTMASK = 16'h5ccf;
    EFX_LUT4 LUT__2844 (.I0(n1642), .I1(n1944), .I2(n703), .O(n1960)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__2844.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__2845 (.I0(n762), .I1(n701), .I2(n1960), .I3(n1646), 
            .O(n1961)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc355 */ ;
    defparam LUT__2845.LUTMASK = 16'hc355;
    EFX_LUT4 LUT__2846 (.I0(n1961), .I1(n1708), .I2(n1959), .I3(n1711), 
            .O(n1962)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__2846.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__2847 (.I0(n1656), .I1(n641), .I2(n1665), .I3(\CPU/cycles[9] ), 
            .O(n1963)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2847.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2848 (.I0(n1957), .I1(n1958), .I2(n1962), .I3(n1963), 
            .O(n1964)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__2848.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__2849 (.I0(n1940), .I1(n1955), .I2(n1954), .I3(n1964), 
            .O(\CPU/writeBackData[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h01ff */ ;
    defparam LUT__2849.LUTMASK = 16'h01ff;
    EFX_LUT4 LUT__2850 (.I0(\mem_rdata[10] ), .I1(\mem_rdata[26] ), .I2(n1611), 
            .I3(n1825), .O(n1965)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__2850.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__2851 (.I0(\CPU/instr[30] ), .I1(\CPU/rs2[10] ), .I2(\CPU/instr[4]~FF_frt_1_frt_2_q ), 
            .O(n1567)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__2851.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__2852 (.I0(\CPU/instr[13] ), .I1(\CPU/instr[12] ), .I2(n1567), 
            .I3(\CPU/rs1[10] ), .O(n1966)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ccf */ ;
    defparam LUT__2852.LUTMASK = 16'h5ccf;
    EFX_LUT4 LUT__2853 (.I0(n1658), .I1(n1948), .I2(\CPU/PC[8] ), .I3(\CPU/PC[9] ), 
            .O(n1967)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2853.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2854 (.I0(n1967), .I1(\CPU/PC[10] ), .O(n1968)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__2854.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__2855 (.I0(n1664), .I1(n1968), .O(n1969)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__2855.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__2856 (.I0(n1656), .I1(n639), .I2(n1665), .I3(\CPU/cycles[10] ), 
            .O(n1970)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2856.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2857 (.I0(n1711), .I1(n1966), .I2(n1969), .I3(n1970), 
            .O(n1971)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__2857.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__2858 (.I0(n1641), .I1(n1642), .I2(n1732), .O(n1972)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__2858.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__2859 (.I0(n760), .I1(n699), .I2(n1972), .I3(n1646), 
            .O(n1973)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc355 */ ;
    defparam LUT__2859.LUTMASK = 16'hc355;
    EFX_LUT4 LUT__2860 (.I0(n1973), .I1(n1708), .I2(\CPU/aluReg[10] ), 
            .I3(n1595), .O(n1974)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bbb */ ;
    defparam LUT__2860.LUTMASK = 16'h0bbb;
    EFX_LUT4 LUT__2861 (.I0(n1965), .I1(n1940), .I2(n1971), .I3(n1974), 
            .O(\CPU/writeBackData[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1fff */ ;
    defparam LUT__2861.LUTMASK = 16'h1fff;
    EFX_LUT4 LUT__2862 (.I0(\mem_rdata[11] ), .I1(\mem_rdata[27] ), .I2(n1611), 
            .I3(n1825), .O(n1975)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__2862.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__2863 (.I0(n1972), .I1(n699), .I2(n697), .I3(n1646), 
            .O(n1976)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8700 */ ;
    defparam LUT__2863.LUTMASK = 16'h8700;
    EFX_LUT4 LUT__2864 (.I0(n758), .I1(n1646), .I2(n1670), .O(n1977)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__2864.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__2865 (.I0(\CPU/rs2[11] ), .I1(\CPU/instr[31] ), .I2(\CPU/instr[4]~FF_frt_1_q ), 
            .I3(\CPU/instr[2]~FF_frt_0_q ), .O(n1565)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__2865.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__2866 (.I0(\CPU/instr[13] ), .I1(\CPU/instr[12] ), .I2(n1565), 
            .I3(\CPU/rs1[11] ), .O(n1978)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ccf */ ;
    defparam LUT__2866.LUTMASK = 16'h5ccf;
    EFX_LUT4 LUT__2867 (.I0(n1594), .I1(\CPU/aluReg[11] ), .I2(n1978), 
            .I3(\CPU/instr[14] ), .O(n1979)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077 */ ;
    defparam LUT__2867.LUTMASK = 16'h7077;
    EFX_LUT4 LUT__2868 (.I0(n1976), .I1(n1977), .I2(n1979), .I3(n1593), 
            .O(n1980)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__2868.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__2869 (.I0(n1967), .I1(\CPU/PC[10] ), .O(n1981)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2869.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2870 (.I0(n1981), .I1(\CPU/PC[11] ), .O(n1982)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__2870.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__2871 (.I0(n1656), .I1(n637), .I2(n1665), .I3(\CPU/cycles[11] ), 
            .O(n1983)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2871.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2872 (.I0(n1664), .I1(n1982), .I2(n1983), .O(n1984)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__2872.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__2873 (.I0(n1975), .I1(n1940), .I2(n1980), .I3(n1984), 
            .O(\CPU/writeBackData[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf1ff */ ;
    defparam LUT__2873.LUTMASK = 16'hf1ff;
    EFX_LUT4 LUT__2874 (.I0(\mem_rdata[12] ), .I1(\mem_rdata[28] ), .I2(n1611), 
            .I3(n1825), .O(n1985)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__2874.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__2875 (.I0(n697), .I1(n699), .O(n1986)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2875.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2876 (.I0(n1641), .I1(n1642), .I2(n1986), .I3(n1732), 
            .O(n1987)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2876.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2877 (.I0(n756), .I1(n695), .I2(n1987), .I3(n1646), 
            .O(n1988)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc355 */ ;
    defparam LUT__2877.LUTMASK = 16'hc355;
    EFX_LUT4 LUT__2878 (.I0(\CPU/rs2[12] ), .I1(\CPU/instr[31] ), .I2(\CPU/instr[4]~FF_frt_1_q ), 
            .I3(\CPU/instr[2]~FF_frt_0_q ), .O(n1563)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__2878.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__2879 (.I0(\CPU/instr[13] ), .I1(\CPU/instr[12] ), .I2(n1563), 
            .I3(\CPU/rs1[12] ), .O(n1989)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ccf */ ;
    defparam LUT__2879.LUTMASK = 16'h5ccf;
    EFX_LUT4 LUT__2880 (.I0(n1594), .I1(\CPU/aluReg[12] ), .I2(n1989), 
            .I3(\CPU/instr[14] ), .O(n1990)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077 */ ;
    defparam LUT__2880.LUTMASK = 16'h7077;
    EFX_LUT4 LUT__2881 (.I0(n1988), .I1(n1670), .I2(n1990), .I3(n1593), 
            .O(n1991)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__2881.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__2882 (.I0(n1981), .I1(\CPU/PC[11] ), .I2(n1664), .I3(\CPU/PC[12] ), 
            .O(n1992)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0708 */ ;
    defparam LUT__2882.LUTMASK = 16'h0708;
    EFX_LUT4 LUT__2883 (.I0(n1656), .I1(n635), .I2(n1665), .I3(\CPU/cycles[12] ), 
            .O(n1993)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2883.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2884 (.I0(\CPU/instr[12] ), .I1(n1666), .I2(n1992), 
            .I3(n1993), .O(n1994)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__2884.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__2885 (.I0(n1985), .I1(n1940), .I2(n1991), .I3(n1994), 
            .O(\CPU/writeBackData[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf1ff */ ;
    defparam LUT__2885.LUTMASK = 16'hf1ff;
    EFX_LUT4 LUT__2886 (.I0(\mem_rdata[13] ), .I1(\mem_rdata[29] ), .I2(n1611), 
            .I3(n1825), .O(n1995)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__2886.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__2887 (.I0(\CPU/instr[31] ), .I1(\CPU/rs2[13] ), .I2(\CPU/instr[4]~FF_frt_1_frt_2_q ), 
            .O(n1561)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__2887.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__2888 (.I0(\CPU/instr[13] ), .I1(\CPU/instr[12] ), .I2(n1561), 
            .I3(\CPU/rs1[13] ), .O(n1996)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ccf */ ;
    defparam LUT__2888.LUTMASK = 16'h5ccf;
    EFX_LUT4 LUT__2889 (.I0(n1987), .I1(n695), .I2(n693), .I3(n1646), 
            .O(n1997)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8700 */ ;
    defparam LUT__2889.LUTMASK = 16'h8700;
    EFX_LUT4 LUT__2890 (.I0(n754), .I1(n1646), .I2(n1997), .I3(n1708), 
            .O(n1998)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__2890.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__2891 (.I0(n1967), .I1(\CPU/PC[10] ), .I2(\CPU/PC[11] ), 
            .I3(\CPU/PC[12] ), .O(n1999)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2891.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2892 (.I0(n633), .I1(\CPU/instr[13] ), .I2(\CPU/instr[5] ), 
            .I3(n1655), .O(n2000)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__2892.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__2893 (.I0(\CPU/instr[2]~FF_frt_0_q ), .I1(\CPU/instr[4] ), 
            .I2(\CPU/instr[6] ), .I3(\CPU/cycles[13] ), .O(n2001)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2893.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2894 (.I0(n1593), .I1(n1594), .I2(\CPU/aluReg[13] ), 
            .O(n2002)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__2894.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__2895 (.I0(n1654), .I1(n2000), .I2(n2001), .I3(n2002), 
            .O(n2003)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__2895.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__2896 (.I0(n1664), .I1(n1999), .I2(\CPU/PC[13] ), .I3(n2003), 
            .O(n2004)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb00 */ ;
    defparam LUT__2896.LUTMASK = 16'heb00;
    EFX_LUT4 LUT__2897 (.I0(n1711), .I1(n1996), .I2(n1998), .I3(n2004), 
            .O(n2005)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__2897.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__2898 (.I0(n1995), .I1(n1940), .I2(n2005), .O(\CPU/writeBackData[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f1f */ ;
    defparam LUT__2898.LUTMASK = 16'h1f1f;
    EFX_LUT4 LUT__2899 (.I0(n752), .I1(n691), .I2(n1733), .I3(n1646), 
            .O(n2006)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc355 */ ;
    defparam LUT__2899.LUTMASK = 16'hc355;
    EFX_LUT4 LUT__2900 (.I0(\CPU/instr[31] ), .I1(\CPU/rs2[14] ), .I2(\CPU/instr[4]~FF_frt_1_frt_2_q ), 
            .O(n1559)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__2900.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__2901 (.I0(\CPU/instr[13] ), .I1(\CPU/instr[12] ), .I2(n1559), 
            .I3(\CPU/rs1[14] ), .O(n2007)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ccf */ ;
    defparam LUT__2901.LUTMASK = 16'h5ccf;
    EFX_LUT4 LUT__2902 (.I0(n2007), .I1(n1711), .I2(n2006), .I3(n1708), 
            .O(n2008)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__2902.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__2903 (.I0(\mem_rdata[14] ), .I1(\mem_rdata[30] ), .I2(n1611), 
            .I3(n1825), .O(n2009)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__2903.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__2904 (.I0(n1661), .I1(\CPU/PC[14] ), .O(n2010)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__2904.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__2905 (.I0(n631), .I1(\CPU/instr[14] ), .I2(\CPU/instr[5] ), 
            .I3(n1655), .O(n2011)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__2905.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__2906 (.I0(\CPU/instr[2]~FF_frt_0_q ), .I1(\CPU/instr[4] ), 
            .I2(\CPU/instr[6] ), .I3(\CPU/cycles[14] ), .O(n2012)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2906.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2907 (.I0(n1593), .I1(n1594), .I2(\CPU/aluReg[14] ), 
            .O(n2013)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__2907.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__2908 (.I0(n1654), .I1(n2011), .I2(n2012), .I3(n2013), 
            .O(n2014)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__2908.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__2909 (.I0(n1664), .I1(n2010), .I2(n2014), .O(n2015)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__2909.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__2910 (.I0(n2009), .I1(n1940), .I2(n2008), .I3(n2015), 
            .O(\CPU/writeBackData[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1fff */ ;
    defparam LUT__2910.LUTMASK = 16'h1fff;
    EFX_LUT4 LUT__2911 (.I0(n1633), .I1(\mem_rdata[15] ), .I2(\CPU/instr[13] ), 
            .O(n2016)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__2911.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__2912 (.I0(n1643), .I1(n691), .I2(n701), .O(n2017)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__2912.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__2913 (.I0(n1960), .I1(n2017), .I2(n689), .I3(n1646), 
            .O(n2018)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8700 */ ;
    defparam LUT__2913.LUTMASK = 16'h8700;
    EFX_LUT4 LUT__2914 (.I0(n750), .I1(n1646), .I2(n2018), .I3(n1708), 
            .O(n2019)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__2914.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__2915 (.I0(n1661), .I1(\CPU/PC[14] ), .I2(n1664), .I3(\CPU/PC[15] ), 
            .O(n2020)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0708 */ ;
    defparam LUT__2915.LUTMASK = 16'h0708;
    EFX_LUT4 LUT__2916 (.I0(\CPU/rs2[15] ), .I1(\CPU/instr[31] ), .I2(\CPU/instr[4]~FF_frt_1_q ), 
            .I3(\CPU/instr[2]~FF_frt_0_q ), .O(n1557)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc */ ;
    defparam LUT__2916.LUTMASK = 16'haccc;
    EFX_LUT4 LUT__2917 (.I0(\CPU/instr[13] ), .I1(\CPU/instr[12] ), .I2(n1557), 
            .I3(\CPU/rs1[15] ), .O(n2021)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ccf */ ;
    defparam LUT__2917.LUTMASK = 16'h5ccf;
    EFX_LUT4 LUT__2918 (.I0(\CPU/instr[15] ), .I1(n1666), .I2(n1665), 
            .I3(\CPU/cycles[15] ), .O(n2022)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2918.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2919 (.I0(n1656), .I1(n629), .I2(n1595), .I3(\CPU/aluReg[15] ), 
            .O(n2023)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__2919.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__2920 (.I0(n1711), .I1(n2021), .I2(n2022), .I3(n2023), 
            .O(n2024)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd000 */ ;
    defparam LUT__2920.LUTMASK = 16'hd000;
    EFX_LUT4 LUT__2921 (.I0(n2019), .I1(n2020), .I2(n2024), .O(n2025)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__2921.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__2922 (.I0(n1940), .I1(n2016), .I2(n2025), .O(\CPU/writeBackData[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f1f */ ;
    defparam LUT__2922.LUTMASK = 16'h1f1f;
    EFX_LUT4 LUT__2923 (.I0(\CPU/instr[14] ), .I1(n1594), .O(n2026)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__2923.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__2924 (.I0(\CPU/aluReg[2] ), .I1(\CPU/aluReg[0] ), .I2(n2026), 
            .O(n2027)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__2924.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__2925 (.I0(n2027), .I1(\CPU/rs1[1] ), .I2(n1592), .O(\CPU/n1066 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__2925.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__2926 (.I0(n2026), .I1(\CPU/aluReg[1] ), .I2(\CPU/rs1[0] ), 
            .I3(n1592), .O(\CPU/n1067 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044 */ ;
    defparam LUT__2926.LUTMASK = 16'hf044;
    EFX_LUT4 LUT__2927 (.I0(n1585), .I1(n1592), .I2(\CPU/aluShamt[0] ), 
            .I3(\CPU/aluShamt[1] ), .O(\CPU/n1033 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb00b */ ;
    defparam LUT__2927.LUTMASK = 16'hb00b;
    EFX_LUT4 LUT__2928 (.I0(\CPU/aluShamt[0] ), .I1(\CPU/aluShamt[1] ), 
            .I2(\CPU/aluShamt[2] ), .O(n2028)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he1e1 */ ;
    defparam LUT__2928.LUTMASK = 16'he1e1;
    EFX_LUT4 LUT__2929 (.I0(n1583), .I1(n1592), .I2(n2028), .O(\CPU/n1032 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__2929.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__2930 (.I0(\CPU/aluShamt[4] ), .I1(n1581), .I2(\CPU/aluShamt[3] ), 
            .I3(n1590), .O(\CPU/n1031 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0ef0 */ ;
    defparam LUT__2930.LUTMASK = 16'h0ef0;
    EFX_LUT4 LUT__2931 (.I0(n1579), .I1(\CPU/aluShamt[4] ), .I2(n1591), 
            .O(\CPU/n1030 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2c2c */ ;
    defparam LUT__2931.LUTMASK = 16'h2c2c;
    EFX_LUT4 LUT__2932 (.I0(\CPU/state[2] ), .I1(n1592), .I2(\CPU/state[1] ), 
            .I3(\CPU/state[3] ), .O(\CPU/select_174/Select_1/n5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3005 */ ;
    defparam LUT__2932.LUTMASK = 16'h3005;
    EFX_LUT4 LUT__2933 (.I0(n1592), .I1(\CPU/state[2] ), .I2(\CPU/state[3] ), 
            .I3(\CPU/state[1] ), .O(\CPU/n2183 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40 */ ;
    defparam LUT__2933.LUTMASK = 16'hff40;
    EFX_LUT4 LUT__2934 (.I0(\CPU/state[2] ), .I1(n1597), .I2(n1592), .I3(\CPU/state[3] ), 
            .O(\CPU/n2182 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f88 */ ;
    defparam LUT__2934.LUTMASK = 16'h8f88;
    EFX_LUT4 LUT__2935 (.I0(n1663), .I1(n1654), .O(n2029)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2935.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2936 (.I0(n8), .I1(n778), .I2(n2029), .O(\CPU/n2063 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__2936.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__2937 (.I0(n1645), .I1(n1835), .I2(\CPU/instr[12] ), 
            .O(n2030)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8787 */ ;
    defparam LUT__2937.LUTMASK = 16'h8787;
    EFX_LUT4 LUT__2938 (.I0(n658), .I1(\CPU/instr[14] ), .I2(\CPU/instr[13] ), 
            .O(n2031)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7c7c */ ;
    defparam LUT__2938.LUTMASK = 16'h7c7c;
    EFX_LUT4 LUT__2939 (.I0(n1596), .I1(n1663), .O(n2032)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2939.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2940 (.I0(n1649), .I1(n2030), .I2(n2031), .I3(n2032), 
            .O(n2033)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8300 */ ;
    defparam LUT__2940.LUTMASK = 16'h8300;
    EFX_LUT4 LUT__2941 (.I0(n2032), .I1(n1594), .I2(\CPU/instr[14] ), 
            .O(n2034)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__2941.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__2942 (.I0(\CPU/rs1[31] ), .I1(n1836), .I2(n1525), .I3(n2034), 
            .O(n2035)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd000 */ ;
    defparam LUT__2942.LUTMASK = 16'hd000;
    EFX_LUT4 LUT__2943 (.I0(\CPU/rs1[31] ), .I1(n1594), .I2(n2032), .I3(\CPU/instr[14] ), 
            .O(n2036)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__2943.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__2944 (.I0(n1596), .I1(n1611), .I2(n1663), .I3(\CPU/instr[14] ), 
            .O(n2037)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__2944.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__2945 (.I0(\CPU/rs1[31] ), .I1(n1525), .I2(n2037), .O(n2038)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__2945.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__2946 (.I0(n1525), .I1(n2037), .I2(\CPU/rs1[31] ), .I3(\CPU/instr[3] ), 
            .O(n2039)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf */ ;
    defparam LUT__2946.LUTMASK = 16'h00bf;
    EFX_LUT4 LUT__2947 (.I0(n2038), .I1(n2036), .I2(n1836), .I3(n2039), 
            .O(n2040)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__2947.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__2948 (.I0(n2033), .I1(n2035), .I2(n2040), .O(n2041)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__2948.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__2949 (.I0(n2041), .I1(n1664), .I2(resetn), .I3(\CPU/state[2] ), 
            .O(ceg_net32)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00 */ ;
    defparam LUT__2949.LUTMASK = 16'h7f00;
    EFX_LUT4 LUT__2950 (.I0(n2035), .I1(n2033), .I2(n2040), .I3(n655), 
            .O(n2042)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__2950.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__2951 (.I0(n2033), .I1(n2035), .I2(\CPU/PC[2] ), .I3(n2040), 
            .O(n2043)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__2951.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__2952 (.I0(n2043), .I1(n2042), .I2(n776), .I3(n2029), 
            .O(\CPU/n2062 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__2952.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__2953 (.I0(n2035), .I1(n2033), .I2(n2040), .I3(n653), 
            .O(n2044)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__2953.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__2954 (.I0(n2033), .I1(n2035), .I2(n1884), .I3(n2040), 
            .O(n2045)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__2954.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__2955 (.I0(n2045), .I1(n2044), .I2(n774), .I3(n2029), 
            .O(\CPU/n2061 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011 */ ;
    defparam LUT__2955.LUTMASK = 16'hf011;
    EFX_LUT4 LUT__2956 (.I0(n2035), .I1(n2033), .I2(n2040), .I3(n651), 
            .O(n2046)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__2956.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__2957 (.I0(n2033), .I1(n2035), .I2(n1891), .I3(n2040), 
            .O(n2047)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__2957.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__2958 (.I0(n2047), .I1(n2046), .I2(n772), .I3(n2029), 
            .O(\CPU/n2060 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011 */ ;
    defparam LUT__2958.LUTMASK = 16'hf011;
    EFX_LUT4 LUT__2959 (.I0(n2035), .I1(n2033), .I2(n2040), .I3(n649), 
            .O(n2048)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__2959.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__2960 (.I0(n2033), .I1(n2035), .I2(n1903), .I3(n2040), 
            .O(n2049)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__2960.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__2961 (.I0(n2049), .I1(n2048), .I2(n770), .I3(n2029), 
            .O(\CPU/n2059 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011 */ ;
    defparam LUT__2961.LUTMASK = 16'hf011;
    EFX_LUT4 LUT__2962 (.I0(n2035), .I1(n2033), .I2(n2040), .I3(n647), 
            .O(n2050)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__2962.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__2963 (.I0(n2033), .I1(n2035), .I2(n1922), .I3(n2040), 
            .O(n2051)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__2963.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__2964 (.I0(n2051), .I1(n2050), .I2(n768), .I3(n2029), 
            .O(\CPU/n2058 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011 */ ;
    defparam LUT__2964.LUTMASK = 16'hf011;
    EFX_LUT4 LUT__2965 (.I0(n2035), .I1(n2033), .I2(n2040), .I3(n645), 
            .O(n2052)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__2965.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__2966 (.I0(n2033), .I1(n2035), .I2(n1934), .I3(n2040), 
            .O(n2053)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__2966.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__2967 (.I0(n2053), .I1(n2052), .I2(n766), .I3(n2029), 
            .O(\CPU/n2057 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011 */ ;
    defparam LUT__2967.LUTMASK = 16'hf011;
    EFX_LUT4 LUT__2968 (.I0(n2035), .I1(n2033), .I2(n2040), .I3(n643), 
            .O(n2054)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__2968.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__2969 (.I0(n2033), .I1(n2035), .I2(n1950), .I3(n2040), 
            .O(n2055)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__2969.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__2970 (.I0(n2055), .I1(n2054), .I2(n764), .I3(n2029), 
            .O(\CPU/n2056 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011 */ ;
    defparam LUT__2970.LUTMASK = 16'hf011;
    EFX_LUT4 LUT__2971 (.I0(n2035), .I1(n2033), .I2(n2040), .I3(n641), 
            .O(n2056)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__2971.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__2972 (.I0(n2033), .I1(n2035), .I2(n1956), .I3(n2040), 
            .O(n2057)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__2972.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__2973 (.I0(n2057), .I1(n2056), .I2(n762), .I3(n2029), 
            .O(\CPU/n2055 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011 */ ;
    defparam LUT__2973.LUTMASK = 16'hf011;
    EFX_LUT4 LUT__2974 (.I0(n2035), .I1(n2033), .I2(n2040), .I3(n639), 
            .O(n2058)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__2974.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__2975 (.I0(n2033), .I1(n2035), .I2(n1968), .I3(n2040), 
            .O(n2059)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__2975.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__2976 (.I0(n2059), .I1(n2058), .I2(n760), .I3(n2029), 
            .O(\CPU/n2054 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011 */ ;
    defparam LUT__2976.LUTMASK = 16'hf011;
    EFX_LUT4 LUT__2977 (.I0(n2035), .I1(n2033), .I2(n2040), .I3(n637), 
            .O(n2060)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__2977.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__2978 (.I0(n2033), .I1(n2035), .I2(n1982), .I3(n2040), 
            .O(n2061)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__2978.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__2979 (.I0(n2061), .I1(n2060), .I2(n758), .I3(n2029), 
            .O(\CPU/n2053 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011 */ ;
    defparam LUT__2979.LUTMASK = 16'hf011;
    EFX_LUT4 LUT__2980 (.I0(n1981), .I1(\CPU/PC[11] ), .I2(\CPU/PC[12] ), 
            .O(n2062)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__2980.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__2981 (.I0(n2033), .I1(n2035), .I2(n2062), .I3(n2040), 
            .O(n2063)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__2981.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__2982 (.I0(n2035), .I1(n2033), .I2(n2040), .I3(n635), 
            .O(n2064)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__2982.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__2983 (.I0(n2064), .I1(n2063), .I2(n756), .I3(n2029), 
            .O(\CPU/n2052 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011 */ ;
    defparam LUT__2983.LUTMASK = 16'hf011;
    EFX_LUT4 LUT__2984 (.I0(n2035), .I1(n2033), .I2(n2040), .I3(n633), 
            .O(n2065)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__2984.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__2985 (.I0(n1999), .I1(\CPU/PC[13] ), .O(n2066)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__2985.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__2986 (.I0(n2033), .I1(n2035), .I2(n2066), .I3(n2040), 
            .O(n2067)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__2986.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__2987 (.I0(n2067), .I1(n2065), .I2(n754), .I3(n2029), 
            .O(\CPU/n2051 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011 */ ;
    defparam LUT__2987.LUTMASK = 16'hf011;
    EFX_LUT4 LUT__2988 (.I0(n2035), .I1(n2033), .I2(n2040), .I3(n631), 
            .O(n2068)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__2988.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__2989 (.I0(n2033), .I1(n2035), .I2(n2010), .I3(n2040), 
            .O(n2069)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__2989.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__2990 (.I0(n2069), .I1(n2068), .I2(n752), .I3(n2029), 
            .O(\CPU/n2050 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011 */ ;
    defparam LUT__2990.LUTMASK = 16'hf011;
    EFX_LUT4 LUT__2991 (.I0(n1661), .I1(\CPU/PC[14] ), .I2(n2029), .I3(\CPU/PC[15] ), 
            .O(n2070)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0708 */ ;
    defparam LUT__2991.LUTMASK = 16'h0708;
    EFX_LUT4 LUT__2992 (.I0(n2029), .I1(n750), .O(n2071)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__2992.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__2993 (.I0(n629), .I1(n2070), .I2(n2071), .I3(n2041), 
            .O(\CPU/n2049 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfcfa */ ;
    defparam LUT__2993.LUTMASK = 16'hfcfa;
    EFX_LUT4 LUT__2994 (.I0(n2033), .I1(n2035), .I2(n1662), .I3(n2040), 
            .O(n2072)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__2994.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__2995 (.I0(n2035), .I1(n2033), .I2(n2040), .I3(n627), 
            .O(n2073)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__2995.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__2996 (.I0(n2073), .I1(n2072), .I2(n748), .I3(n2029), 
            .O(\CPU/n2048 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011 */ ;
    defparam LUT__2996.LUTMASK = 16'hf011;
    EFX_LUT4 LUT__2997 (.I0(n2035), .I1(n2033), .I2(n2040), .I3(n625), 
            .O(n2074)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__2997.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__2998 (.I0(n1661), .I1(n1677), .I2(\CPU/PC[17] ), .O(n2075)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__2998.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__2999 (.I0(n2033), .I1(n2035), .I2(n2075), .I3(n2040), 
            .O(n2076)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__2999.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__3000 (.I0(n2076), .I1(n2074), .I2(n746), .I3(n2029), 
            .O(\CPU/n2047 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011 */ ;
    defparam LUT__3000.LUTMASK = 16'hf011;
    EFX_LUT4 LUT__3001 (.I0(n2035), .I1(n2033), .I2(n2040), .I3(n623), 
            .O(n2077)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__3001.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__3002 (.I0(n1689), .I1(\CPU/PC[18] ), .O(n2078)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3002.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3003 (.I0(n2033), .I1(n2035), .I2(n2078), .I3(n2040), 
            .O(n2079)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__3003.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__3004 (.I0(n2079), .I1(n2077), .I2(n744), .I3(n2029), 
            .O(\CPU/n2046 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011 */ ;
    defparam LUT__3004.LUTMASK = 16'hf011;
    EFX_LUT4 LUT__3005 (.I0(n2035), .I1(n2033), .I2(n2040), .I3(n621), 
            .O(n2080)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__3005.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__3006 (.I0(n1699), .I1(\CPU/PC[19] ), .O(n2081)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3006.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3007 (.I0(n2033), .I1(n2035), .I2(n2081), .I3(n2040), 
            .O(n2082)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__3007.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__3008 (.I0(n2082), .I1(n2080), .I2(n742), .I3(n2029), 
            .O(\CPU/n2045 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011 */ ;
    defparam LUT__3008.LUTMASK = 16'hf011;
    EFX_LUT4 LUT__3009 (.I0(n2035), .I1(n2033), .I2(n2040), .I3(n619), 
            .O(n2083)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__3009.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__3010 (.I0(n2033), .I1(n2035), .I2(n1704), .I3(n2040), 
            .O(n2084)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__3010.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__3011 (.I0(n2084), .I1(n2083), .I2(n740), .I3(n2029), 
            .O(\CPU/n2044 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011 */ ;
    defparam LUT__3011.LUTMASK = 16'hf011;
    EFX_LUT4 LUT__3012 (.I0(n2035), .I1(n2033), .I2(n2040), .I3(n617), 
            .O(n2085)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__3012.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__3013 (.I0(n1699), .I1(n1723), .I2(\CPU/PC[21] ), .O(n2086)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__3013.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__3014 (.I0(n2033), .I1(n2035), .I2(n2086), .I3(n2040), 
            .O(n2087)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__3014.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__3015 (.I0(n2087), .I1(n2085), .I2(n738), .I3(n2029), 
            .O(\CPU/n2043 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011 */ ;
    defparam LUT__3015.LUTMASK = 16'hf011;
    EFX_LUT4 LUT__3016 (.I0(n2035), .I1(n2033), .I2(n2040), .I3(n615), 
            .O(n2088)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__3016.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__3017 (.I0(n2033), .I1(n2035), .I2(n1728), .I3(n2040), 
            .O(n2089)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__3017.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__3018 (.I0(n2089), .I1(n2088), .I2(n736), .I3(n2029), 
            .O(\CPU/n2042 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011 */ ;
    defparam LUT__3018.LUTMASK = 16'hf011;
    EFX_LUT4 LUT__3019 (.I0(n2033), .I1(n2035), .I2(n1743), .I3(n2040), 
            .O(n2090)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__3019.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__3020 (.I0(n2035), .I1(n2033), .I2(n2040), .I3(n614), 
            .O(n2091)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__3020.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__3021 (.I0(n2091), .I1(n2090), .I2(n734), .I3(n2029), 
            .O(\CPU/n2041 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011 */ ;
    defparam LUT__3021.LUTMASK = 16'hf011;
    EFX_LUT4 LUT__3022 (.I0(\CPU/aluReg[3] ), .I1(\CPU/aluReg[1] ), .I2(n2026), 
            .O(n2092)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3022.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3023 (.I0(n2092), .I1(\CPU/rs1[2] ), .I2(n1592), .O(\CPU/n1065 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__3023.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__3024 (.I0(\CPU/aluReg[4] ), .I1(\CPU/aluReg[2] ), .I2(n2026), 
            .O(n2093)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3024.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3025 (.I0(n2093), .I1(\CPU/rs1[3] ), .I2(n1592), .O(\CPU/n1064 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__3025.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__3026 (.I0(\CPU/aluReg[5] ), .I1(\CPU/aluReg[3] ), .I2(n2026), 
            .O(n2094)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3026.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3027 (.I0(n2094), .I1(\CPU/rs1[4] ), .I2(n1592), .O(\CPU/n1063 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__3027.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__3028 (.I0(\CPU/aluReg[6] ), .I1(\CPU/aluReg[4] ), .I2(n2026), 
            .O(n2095)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3028.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3029 (.I0(n2095), .I1(\CPU/rs1[5] ), .I2(n1592), .O(\CPU/n1062 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__3029.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__3030 (.I0(\CPU/aluReg[7] ), .I1(\CPU/aluReg[5] ), .I2(n2026), 
            .O(n2096)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3030.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3031 (.I0(n2096), .I1(\CPU/rs1[6] ), .I2(n1592), .O(\CPU/n1061 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__3031.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__3032 (.I0(\CPU/aluReg[8] ), .I1(\CPU/aluReg[6] ), .I2(n2026), 
            .O(n2097)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3032.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3033 (.I0(n2097), .I1(\CPU/rs1[7] ), .I2(n1592), .O(\CPU/n1060 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__3033.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__3034 (.I0(\CPU/aluReg[9] ), .I1(\CPU/aluReg[7] ), .I2(n2026), 
            .O(n2098)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3034.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3035 (.I0(n2098), .I1(\CPU/rs1[8] ), .I2(n1592), .O(\CPU/n1059 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__3035.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__3036 (.I0(\CPU/aluReg[10] ), .I1(\CPU/aluReg[8] ), .I2(n2026), 
            .O(n2099)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3036.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3037 (.I0(n2099), .I1(\CPU/rs1[9] ), .I2(n1592), .O(\CPU/n1058 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__3037.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__3038 (.I0(\CPU/aluReg[11] ), .I1(\CPU/aluReg[9] ), .I2(n2026), 
            .O(n2100)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3038.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3039 (.I0(n2100), .I1(\CPU/rs1[10] ), .I2(n1592), .O(\CPU/n1057 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3039.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3040 (.I0(\CPU/aluReg[12] ), .I1(\CPU/aluReg[10] ), .I2(n2026), 
            .O(n2101)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3040.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3041 (.I0(n2101), .I1(\CPU/rs1[11] ), .I2(n1592), .O(\CPU/n1056 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3041.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3042 (.I0(\CPU/aluReg[13] ), .I1(\CPU/aluReg[11] ), .I2(n2026), 
            .O(n2102)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3042.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3043 (.I0(n2102), .I1(\CPU/rs1[12] ), .I2(n1592), .O(\CPU/n1055 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__3043.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__3044 (.I0(\CPU/aluReg[14] ), .I1(\CPU/aluReg[12] ), .I2(n2026), 
            .O(n2103)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3044.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3045 (.I0(n2103), .I1(\CPU/rs1[13] ), .I2(n1592), .O(\CPU/n1054 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__3045.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__3046 (.I0(\CPU/aluReg[15] ), .I1(\CPU/aluReg[13] ), .I2(n2026), 
            .O(n2104)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3046.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3047 (.I0(n2104), .I1(\CPU/rs1[14] ), .I2(n1592), .O(\CPU/n1053 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3047.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3048 (.I0(\CPU/aluReg[16] ), .I1(\CPU/aluReg[14] ), .I2(n2026), 
            .O(n2105)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3048.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3049 (.I0(n2105), .I1(\CPU/rs1[15] ), .I2(n1592), .O(\CPU/n1052 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3049.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3050 (.I0(\CPU/aluReg[17] ), .I1(\CPU/aluReg[15] ), .I2(n2026), 
            .O(n2106)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3050.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3051 (.I0(n2106), .I1(\CPU/rs1[16] ), .I2(n1592), .O(\CPU/n1051 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3051.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3052 (.I0(\CPU/aluReg[18] ), .I1(\CPU/aluReg[16] ), .I2(n2026), 
            .O(n2107)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3052.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3053 (.I0(n2107), .I1(\CPU/rs1[17] ), .I2(n1592), .O(\CPU/n1050 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__3053.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__3054 (.I0(\CPU/aluReg[19] ), .I1(\CPU/aluReg[17] ), .I2(n2026), 
            .O(n2108)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3054.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3055 (.I0(n2108), .I1(\CPU/rs1[18] ), .I2(n1592), .O(\CPU/n1049 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__3055.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__3056 (.I0(\CPU/aluReg[20] ), .I1(\CPU/aluReg[18] ), .I2(n2026), 
            .O(n2109)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3056.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3057 (.I0(n2109), .I1(\CPU/rs1[19] ), .I2(n1592), .O(\CPU/n1048 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__3057.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__3058 (.I0(\CPU/aluReg[21] ), .I1(\CPU/aluReg[19] ), .I2(n2026), 
            .O(n2110)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3058.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3059 (.I0(n2110), .I1(\CPU/rs1[20] ), .I2(n1592), .O(\CPU/n1047 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__3059.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__3060 (.I0(\CPU/aluReg[22] ), .I1(\CPU/aluReg[20] ), .I2(n2026), 
            .O(n2111)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3060.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3061 (.I0(n2111), .I1(\CPU/rs1[21] ), .I2(n1592), .O(\CPU/n1046 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3061.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3062 (.I0(\CPU/aluReg[23] ), .I1(\CPU/aluReg[21] ), .I2(n2026), 
            .O(n2112)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3062.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3063 (.I0(n2112), .I1(\CPU/rs1[22] ), .I2(n1592), .O(\CPU/n1045 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__3063.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__3064 (.I0(\CPU/aluReg[24] ), .I1(\CPU/aluReg[22] ), .I2(n2026), 
            .O(n2113)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3064.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3065 (.I0(n2113), .I1(\CPU/rs1[23] ), .I2(n1592), .O(\CPU/n1044 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3065.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3066 (.I0(\CPU/aluReg[25] ), .I1(\CPU/aluReg[23] ), .I2(n2026), 
            .O(n2114)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3066.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3067 (.I0(n2114), .I1(\CPU/rs1[24] ), .I2(n1592), .O(\CPU/n1043 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3067.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3068 (.I0(\CPU/aluReg[26] ), .I1(\CPU/aluReg[24] ), .I2(n2026), 
            .O(n2115)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3068.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3069 (.I0(n2115), .I1(\CPU/rs1[25] ), .I2(n1592), .O(\CPU/n1042 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3069.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3070 (.I0(\CPU/aluReg[27] ), .I1(\CPU/aluReg[25] ), .I2(n2026), 
            .O(n2116)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3070.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3071 (.I0(n2116), .I1(\CPU/rs1[26] ), .I2(n1592), .O(\CPU/n1041 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3071.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3072 (.I0(\CPU/aluReg[28] ), .I1(\CPU/aluReg[26] ), .I2(n2026), 
            .O(n2117)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3072.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3073 (.I0(n2117), .I1(\CPU/rs1[27] ), .I2(n1592), .O(\CPU/n1040 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__3073.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__3074 (.I0(\CPU/aluReg[29] ), .I1(\CPU/aluReg[27] ), .I2(n2026), 
            .O(n2118)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3074.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3075 (.I0(n2118), .I1(\CPU/rs1[28] ), .I2(n1592), .O(\CPU/n1039 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3075.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3076 (.I0(\CPU/aluReg[30] ), .I1(\CPU/aluReg[28] ), .I2(n2026), 
            .O(n2119)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3076.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3077 (.I0(n2119), .I1(\CPU/rs1[29] ), .I2(n1592), .O(\CPU/n1038 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3077.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3078 (.I0(\CPU/aluReg[31] ), .I1(\CPU/aluReg[29] ), .I2(n2026), 
            .O(n2120)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3078.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3079 (.I0(n2120), .I1(\CPU/rs1[30] ), .I2(n1592), .O(\CPU/n1037 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3079.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3080 (.I0(\CPU/instr[30] ), .I1(\CPU/aluReg[31] ), .I2(\CPU/aluReg[30] ), 
            .I3(n2026), .O(n2121)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f77 */ ;
    defparam LUT__3080.LUTMASK = 16'h0f77;
    EFX_LUT4 LUT__3081 (.I0(n2121), .I1(\CPU/rs1[31] ), .I2(n1592), .O(\CPU/n1036 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__3081.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__3082 (.I0(n1619), .I1(n1830), .O(\RAM/n104 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3082.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3083 (.I0(\CPU/rs2[16] ), .I1(\mem_wdata[0] ), .I2(n612), 
            .O(\mem_wdata[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3083.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3084 (.I0(n1823), .I1(n1620), .O(\RAM/n112 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3084.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3085 (.I0(\CPU/rs2[9] ), .I1(\mem_wdata[1] ), .I2(n12), 
            .O(\mem_wdata[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3085.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3086 (.I0(\mem_wdata[9] ), .I1(\CPU/rs2[25] ), .I2(n1610), 
            .O(\mem_wdata[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3086.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3087 (.I0(\CPU/rs2[10] ), .I1(\mem_wdata[2] ), .I2(n12), 
            .O(\mem_wdata[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3087.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3088 (.I0(n12), .I1(n1611), .I2(n1825), .I3(n1619), 
            .O(\RAM/n108 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__3088.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__3089 (.I0(\mem_wdata[10] ), .I1(\CPU/rs2[26] ), .I2(n1610), 
            .O(\mem_wdata[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3089.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3090 (.I0(\CPU/rs2[18] ), .I1(\mem_wdata[2] ), .I2(n612), 
            .O(\mem_wdata[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3090.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3091 (.I0(\CPU/rs2[11] ), .I1(\mem_wdata[3] ), .I2(n12), 
            .O(\mem_wdata[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3091.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3092 (.I0(\mem_wdata[11] ), .I1(\CPU/rs2[27] ), .I2(n1610), 
            .O(\mem_wdata[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3092.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3093 (.I0(\CPU/rs2[12] ), .I1(\mem_wdata[4] ), .I2(n12), 
            .O(\mem_wdata[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3093.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3094 (.I0(\mem_wdata[12] ), .I1(\CPU/rs2[28] ), .I2(n1610), 
            .O(\mem_wdata[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3094.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3095 (.I0(\CPU/rs2[13] ), .I1(\mem_wdata[5] ), .I2(n12), 
            .O(\mem_wdata[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3095.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3096 (.I0(\mem_wdata[13] ), .I1(\CPU/rs2[29] ), .I2(n1610), 
            .O(\mem_wdata[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3096.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3097 (.I0(\CPU/rs2[14] ), .I1(\mem_wdata[6] ), .I2(n12), 
            .O(\mem_wdata[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3097.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3098 (.I0(\mem_wdata[14] ), .I1(\CPU/rs2[30] ), .I2(n1610), 
            .O(\mem_wdata[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3098.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3099 (.I0(\CPU/rs2[15] ), .I1(\mem_wdata[7] ), .I2(n12), 
            .O(\mem_wdata[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3099.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3100 (.I0(\mem_wdata[15] ), .I1(\CPU/rs2[31] ), .I2(n1610), 
            .O(\mem_wdata[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3100.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3101 (.I0(\CPU/rs2[17] ), .I1(\mem_wdata[1] ), .I2(n612), 
            .O(\mem_wdata[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3101.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3102 (.I0(\CPU/rs2[19] ), .I1(\mem_wdata[3] ), .I2(n612), 
            .O(\mem_wdata[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3102.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3103 (.I0(\CPU/rs2[20] ), .I1(\mem_wdata[4] ), .I2(n612), 
            .O(\mem_wdata[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3103.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3104 (.I0(\CPU/rs2[21] ), .I1(\mem_wdata[5] ), .I2(n612), 
            .O(\mem_wdata[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3104.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3105 (.I0(\CPU/rs2[22] ), .I1(\mem_wdata[6] ), .I2(n612), 
            .O(\mem_wdata[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3105.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3106 (.I0(\CPU/rs2[23] ), .I1(\mem_wdata[7] ), .I2(n612), 
            .O(\mem_wdata[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3106.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3107 (.I0(\CPU/PC[1] ), .I1(n1610), .I2(n1606), .O(n2122)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__3107.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__3108 (.I0(n2122), .I1(\mem_addr[4] ), .O(n2123)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3108.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3109 (.I0(\mem_addr[2] ), .I1(\mem_addr[3] ), .I2(n1861), 
            .I3(n2123), .O(n2124)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__3109.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__3110 (.I0(n2124), .I1(n1612), .O(\per_uart/n25 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3110.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3111 (.I0(\mem_addr[4] ), .I1(n2122), .O(n2125)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3111.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3112 (.I0(\mem_addr[2] ), .I1(n2125), .I2(n1861), .I3(\mem_addr[3] ), 
            .O(n2126)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__3112.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__3113 (.I0(n2126), .I1(\per_uart/rx_data[0] ), .O(\per_uart/select_21/Select_0/n3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3113.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3114 (.I0(n2126), .I1(n1612), .O(\per_uart/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3114.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3115 (.I0(n2126), .I1(\per_uart/rx_data[1] ), .O(\per_uart/select_21/Select_1/n3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3115.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3116 (.I0(n2126), .I1(\per_uart/rx_data[2] ), .O(\per_uart/select_21/Select_2/n3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3116.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3117 (.I0(n2126), .I1(\per_uart/rx_data[3] ), .O(\per_uart/select_21/Select_3/n3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3117.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3118 (.I0(n2126), .I1(\per_uart/rx_data[4] ), .O(\per_uart/select_21/Select_4/n3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3118.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3119 (.I0(n2126), .I1(\per_uart/rx_data[5] ), .O(\per_uart/select_21/Select_5/n3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3119.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3120 (.I0(n2126), .I1(\per_uart/rx_data[6] ), .O(\per_uart/select_21/Select_6/n3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3120.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3121 (.I0(n2126), .I1(\per_uart/rx_data[7] ), .I2(n2124), 
            .I3(\per_uart/rx_error ), .O(\per_uart/select_21/Select_7/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf888 */ ;
    defparam LUT__3121.LUTMASK = 16'hf888;
    EFX_LUT4 LUT__3122 (.I0(n2124), .I1(\per_uart/rx_avail ), .O(\per_uart/select_21/Select_8/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3122.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3123 (.I0(n2124), .I1(\per_uart/tx_busy ), .O(\per_uart/select_21/Select_9/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3123.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3124 (.I0(\per_uart/uart0/rx_bitcount[1] ), .I1(\per_uart/uart0/rx_bitcount[2] ), 
            .I2(\per_uart/uart0/rx_bitcount[0] ), .I3(\per_uart/uart0/rx_bitcount[3] ), 
            .O(n2127)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1001 */ ;
    defparam LUT__3124.LUTMASK = 16'h1001;
    EFX_LUT4 LUT__3125 (.I0(\per_uart/uart0/rx_bitcount[0] ), .I1(\per_uart/uart0/uart_rxd2 ), 
            .I2(\per_uart/uart0/rx_busy ), .I3(n2127), .O(\per_uart/uart0/n190 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1fff */ ;
    defparam LUT__3125.LUTMASK = 16'h1fff;
    EFX_LUT4 LUT__3126 (.I0(\per_uart/uart0/rx_count16[0] ), .I1(\per_uart/uart0/rx_count16[1] ), 
            .I2(\per_uart/uart0/rx_count16[2] ), .I3(\per_uart/uart0/rx_count16[3] ), 
            .O(n2128)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3126.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3127 (.I0(\per_uart/uart0/uart_rxd2 ), .I1(n2128), .I2(\per_uart/uart0/rx_busy ), 
            .I3(resetn), .O(n2129)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00 */ ;
    defparam LUT__3127.LUTMASK = 16'h3a00;
    EFX_LUT4 LUT__3128 (.I0(\per_uart/uart0/enable16_counter[0] ), .I1(\per_uart/uart0/enable16_counter[1] ), 
            .O(n2130)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__3128.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__3129 (.I0(\per_uart/uart0/enable16_counter[2] ), .I1(\per_uart/uart0/enable16_counter[3] ), 
            .I2(\per_uart/uart0/enable16_counter[4] ), .I3(n2130), .O(n2131)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__3129.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__3130 (.I0(n2129), .I1(n2131), .O(ceg_net530)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3130.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3131 (.I0(\per_uart/uart0/rx_busy ), .I1(\per_uart/uart0/rx_count16[0] ), 
            .O(\per_uart/uart0/n195 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7777 */ ;
    defparam LUT__3131.LUTMASK = 16'h7777;
    EFX_LUT4 LUT__3132 (.I0(\per_uart/uart0/rx_busy ), .I1(\per_uart/uart0/uart_rxd2 ), 
            .I2(resetn), .I3(n2131), .O(ceg_net176)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h40ff */ ;
    defparam LUT__3132.LUTMASK = 16'h40ff;
    EFX_LUT4 LUT__3133 (.I0(\per_uart/uart0/rx_bitcount[0] ), .I1(\per_uart/uart0/rx_busy ), 
            .O(\per_uart/uart0/n200 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3133.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3134 (.I0(n2131), .I1(n2128), .I2(\per_uart/uart0/rx_busy ), 
            .O(n2132)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__3134.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__3135 (.I0(\per_uart/uart0/rx_bitcount[1] ), .I1(\per_uart/uart0/rx_bitcount[2] ), 
            .I2(\per_uart/uart0/rx_bitcount[0] ), .I3(\per_uart/uart0/rx_bitcount[3] ), 
            .O(n2133)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__3135.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__3136 (.I0(n2132), .I1(n2133), .O(n2134)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3136.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3137 (.I0(n2134), .I1(\per_uart/uart0/uart_rxd2 ), .O(\per_uart/uart0/n576 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3137.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3138 (.I0(\per_uart/uart0/n576 ), .I1(resetn), .O(\per_uart/uart0/n581 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3138.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3139 (.I0(\per_uart/uart0/n576 ), .I1(\per_uart/uart_ctrl[1] ), 
            .I2(resetn), .O(ceg_net140)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__3139.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__3140 (.I0(\per_uart/uart0/uart_rxd2 ), .I1(n2134), .O(\per_uart/uart0/n242 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3140.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3141 (.I0(n2134), .I1(\per_uart/uart_ctrl[1] ), .I2(resetn), 
            .O(ceg_net144)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__3141.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__3142 (.I0(n2127), .I1(n2132), .I2(resetn), .O(\per_uart/uart0/n582 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfbf */ ;
    defparam LUT__3142.LUTMASK = 16'hbfbf;
    EFX_LUT4 LUT__3143 (.I0(\per_uart/tx_busy ), .I1(\per_uart/uart_ctrl[0] ), 
            .O(\per_uart/uart0/n316 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3143.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3144 (.I0(\per_uart/uart0/tx_count16[0] ), .I1(n2131), 
            .O(\per_uart/uart0/n422 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3144.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3145 (.I0(\per_uart/uart0/tx_count16[1] ), .I1(\per_uart/uart0/tx_count16[2] ), 
            .I2(\per_uart/uart0/tx_count16[3] ), .I3(\per_uart/tx_busy ), 
            .O(n2135)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__3145.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__3146 (.I0(\per_uart/uart0/n422 ), .I1(n2135), .O(n2136)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3146.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3147 (.I0(\per_uart/uart0/tx_bitcount[2] ), .I1(\per_uart/uart0/tx_bitcount[3] ), 
            .O(n2137)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3147.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3148 (.I0(\per_uart/uart0/tx_bitcount[0] ), .I1(n2137), 
            .I2(\per_uart/uart0/tx_bitcount[1] ), .O(n2138)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3148.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3149 (.I0(n2138), .I1(n2136), .I2(resetn), .O(\per_uart/uart0/n601 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f8f */ ;
    defparam LUT__3149.LUTMASK = 16'h8f8f;
    EFX_LUT4 LUT__3150 (.I0(n2131), .I1(resetn), .O(\per_uart/uart0/n552 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3150.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3151 (.I0(\per_uart/uart0/n552 ), .I1(\per_uart/uart0/n316 ), 
            .O(ceg_net203)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__3151.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__3152 (.I0(\per_uart/uart0/tx_bitcount[2] ), .I1(\per_uart/uart0/tx_bitcount[0] ), 
            .I2(\per_uart/uart0/tx_bitcount[1] ), .I3(\per_uart/uart0/tx_bitcount[3] ), 
            .O(n2139)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1401 */ ;
    defparam LUT__3152.LUTMASK = 16'h1401;
    EFX_LUT4 LUT__3153 (.I0(n2139), .I1(\per_uart/uart0/tx_bitcount[0] ), 
            .I2(\per_uart/uart0/tx_bitcount[3] ), .I3(\per_uart/uart0/txd_reg[0] ), 
            .O(\per_uart/uart0/n386 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfd80 */ ;
    defparam LUT__3153.LUTMASK = 16'hfd80;
    EFX_LUT4 LUT__3154 (.I0(resetn), .I1(n2138), .I2(n2136), .O(ceg_net155)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__3154.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__3155 (.I0(n2139), .I1(n2136), .O(n2140)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3155.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3156 (.I0(\per_uart/d_in_uart[0] ), .I1(\per_uart/uart0/txd_reg[1] ), 
            .I2(n2140), .O(\per_uart/uart0/n438 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3156.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3157 (.I0(\per_uart/uart0/n316 ), .I1(n2140), .I2(resetn), 
            .O(ceg_net159)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__3157.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__3158 (.I0(\per_uart/uart0/tx_bitcount[1] ), .I1(n2137), 
            .I2(\per_uart/uart0/tx_bitcount[0] ), .I3(n2136), .O(\per_uart/uart0/n427 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__3158.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__3159 (.I0(\per_uart/uart0/n316 ), .I1(n2136), .I2(resetn), 
            .O(ceg_net246)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__3159.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__3160 (.I0(\per_uart/uart0/rx_count16[0] ), .I1(\per_uart/uart0/rx_count16[1] ), 
            .I2(\per_uart/uart0/rx_busy ), .O(\per_uart/uart0/n194 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6f6f */ ;
    defparam LUT__3160.LUTMASK = 16'h6f6f;
    EFX_LUT4 LUT__3161 (.I0(\per_uart/uart0/rx_count16[0] ), .I1(\per_uart/uart0/rx_count16[1] ), 
            .I2(\per_uart/uart0/rx_count16[2] ), .I3(\per_uart/uart0/rx_busy ), 
            .O(\per_uart/uart0/n193 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h78ff */ ;
    defparam LUT__3161.LUTMASK = 16'h78ff;
    EFX_LUT4 LUT__3162 (.I0(\per_uart/uart0/rx_count16[0] ), .I1(\per_uart/uart0/rx_count16[1] ), 
            .I2(\per_uart/uart0/rx_count16[2] ), .I3(\per_uart/uart0/rx_count16[3] ), 
            .O(n2141)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__3162.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__3163 (.I0(n2141), .I1(\per_uart/uart0/rx_busy ), .O(\per_uart/uart0/n192 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3163.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3164 (.I0(\per_uart/uart0/rx_bitcount[0] ), .I1(\per_uart/uart0/rx_bitcount[1] ), 
            .I2(\per_uart/uart0/rx_busy ), .O(\per_uart/uart0/n199 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__3164.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__3165 (.I0(\per_uart/uart0/rx_bitcount[0] ), .I1(\per_uart/uart0/rx_bitcount[1] ), 
            .I2(\per_uart/uart0/rx_bitcount[2] ), .I3(\per_uart/uart0/rx_busy ), 
            .O(\per_uart/uart0/n198 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;
    defparam LUT__3165.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__3166 (.I0(\per_uart/uart0/rx_bitcount[0] ), .I1(\per_uart/uart0/rx_bitcount[1] ), 
            .I2(\per_uart/uart0/rx_bitcount[2] ), .I3(\per_uart/uart0/rx_bitcount[3] ), 
            .O(n2142)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__3166.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__3167 (.I0(n2142), .I1(\per_uart/uart0/rx_busy ), .O(\per_uart/uart0/n197 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3167.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3168 (.I0(\per_uart/uart0/tx_count16[0] ), .I1(\per_uart/uart0/tx_count16[1] ), 
            .I2(n2131), .O(\per_uart/uart0/n421 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__3168.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__3169 (.I0(\per_uart/uart0/tx_count16[0] ), .I1(\per_uart/uart0/tx_count16[1] ), 
            .I2(\per_uart/uart0/tx_count16[2] ), .I3(n2131), .O(\per_uart/uart0/n420 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;
    defparam LUT__3169.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__3170 (.I0(\per_uart/uart0/tx_count16[0] ), .I1(\per_uart/uart0/tx_count16[1] ), 
            .I2(\per_uart/uart0/tx_count16[2] ), .I3(\per_uart/uart0/tx_count16[3] ), 
            .O(n2143)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__3170.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__3171 (.I0(n2143), .I1(n2131), .O(\per_uart/uart0/n419 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3171.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3172 (.I0(\per_uart/d_in_uart[1] ), .I1(\per_uart/uart0/txd_reg[2] ), 
            .I2(n2140), .O(\per_uart/uart0/n437 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3172.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3173 (.I0(\per_uart/d_in_uart[2] ), .I1(\per_uart/uart0/txd_reg[3] ), 
            .I2(n2140), .O(\per_uart/uart0/n436 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3173.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3174 (.I0(\per_uart/d_in_uart[3] ), .I1(\per_uart/uart0/txd_reg[4] ), 
            .I2(n2140), .O(\per_uart/uart0/n435 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3174.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3175 (.I0(\per_uart/d_in_uart[4] ), .I1(\per_uart/uart0/txd_reg[5] ), 
            .I2(n2140), .O(\per_uart/uart0/n434 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3175.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3176 (.I0(\per_uart/d_in_uart[5] ), .I1(\per_uart/uart0/txd_reg[6] ), 
            .I2(n2140), .O(\per_uart/uart0/n433 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3176.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3177 (.I0(\per_uart/d_in_uart[6] ), .I1(\per_uart/uart0/txd_reg[7] ), 
            .I2(n2140), .O(\per_uart/uart0/n432 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3177.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3178 (.I0(n2140), .I1(\per_uart/d_in_uart[7] ), .O(\per_uart/uart0/n431 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3178.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3179 (.I0(n2137), .I1(\per_uart/uart0/tx_bitcount[0] ), 
            .I2(\per_uart/uart0/tx_bitcount[1] ), .I3(n2136), .O(\per_uart/uart0/n426 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1c00 */ ;
    defparam LUT__3179.LUTMASK = 16'h1c00;
    EFX_LUT4 LUT__3180 (.I0(\per_uart/uart0/tx_bitcount[0] ), .I1(\per_uart/uart0/tx_bitcount[1] ), 
            .I2(\per_uart/uart0/tx_bitcount[2] ), .I3(n2136), .O(\per_uart/uart0/n425 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;
    defparam LUT__3180.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__3181 (.I0(\per_uart/uart0/tx_bitcount[1] ), .I1(\per_uart/uart0/tx_bitcount[0] ), 
            .I2(\per_uart/uart0/tx_bitcount[2] ), .I3(\per_uart/uart0/tx_bitcount[3] ), 
            .O(n2144)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h827f */ ;
    defparam LUT__3181.LUTMASK = 16'h827f;
    EFX_LUT4 LUT__3182 (.I0(n2144), .I1(n2136), .O(\per_uart/uart0/n424 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3182.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3183 (.I0(\per_uart/uart0/enable16_counter[0] ), .I1(\per_uart/uart0/enable16_counter[1] ), 
            .O(\per_uart/uart0/n732 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__3183.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__3184 (.I0(n2130), .I1(\per_uart/uart0/enable16_counter[2] ), 
            .O(\per_uart/uart0/n737 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3184.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3185 (.I0(\per_uart/uart0/enable16_counter[2] ), .I1(n2130), 
            .I2(\per_uart/uart0/enable16_counter[3] ), .O(\per_uart/uart0/n742 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4 */ ;
    defparam LUT__3185.LUTMASK = 16'hb4b4;
    EFX_LUT4 LUT__3186 (.I0(\per_uart/uart0/enable16_counter[2] ), .I1(\per_uart/uart0/enable16_counter[3] ), 
            .I2(n2130), .I3(\per_uart/uart0/enable16_counter[4] ), .O(\per_uart/uart0/n747 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef10 */ ;
    defparam LUT__3186.LUTMASK = 16'hef10;
    EFX_LUT4 LUT__3187 (.I0(n1622), .I1(n2125), .I2(n1612), .O(n2145)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__3187.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__3188 (.I0(\mem_addr[3] ), .I1(\mem_addr[2] ), .I2(n2145), 
            .O(\mult1/n402 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3188.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3189 (.I0(n2145), .I1(\mem_addr[3] ), .O(n2146)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3189.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3190 (.I0(\mem_addr[2] ), .I1(n2146), .O(\mult1/n403 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3190.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3191 (.I0(\mult1/result[0] ), .I1(\mult1/done ), .I2(\mem_addr[2] ), 
            .O(n2147)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3191.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3192 (.I0(\mem_addr[3] ), .I1(n2123), .I2(n1622), .O(n2148)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3192.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3193 (.I0(\mult_dout[0] ), .I1(n2147), .I2(n2148), .O(\mult1/n201 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3193.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3194 (.I0(n1599), .I1(\CPU/state[2] ), .I2(\CPU/state[0] ), 
            .I3(n1622), .O(\mult1/n165 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__3194.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__3195 (.I0(n2146), .I1(\mem_addr[2] ), .O(\mult1/n404 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3195.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3196 (.I0(\mem_addr[2] ), .I1(\mult1/result[1] ), .I2(\mult_dout[1] ), 
            .I3(n2148), .O(\mult1/n200 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__3196.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__3197 (.I0(\mem_addr[2] ), .I1(\mult1/result[2] ), .I2(\mult_dout[2] ), 
            .I3(n2148), .O(\mult1/n199 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__3197.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__3198 (.I0(\mem_addr[2] ), .I1(\mult1/result[3] ), .I2(\mult_dout[3] ), 
            .I3(n2148), .O(\mult1/n198 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__3198.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__3199 (.I0(\mem_addr[2] ), .I1(\mult1/result[4] ), .I2(\mult_dout[4] ), 
            .I3(n2148), .O(\mult1/n197 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__3199.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__3200 (.I0(\mem_addr[2] ), .I1(\mult1/result[5] ), .I2(\mult_dout[5] ), 
            .I3(n2148), .O(\mult1/n196 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__3200.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__3201 (.I0(\mem_addr[2] ), .I1(\mult1/result[6] ), .I2(\mult_dout[6] ), 
            .I3(n2148), .O(\mult1/n195 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__3201.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__3202 (.I0(\mem_addr[2] ), .I1(\mult1/result[7] ), .I2(\mult_dout[7] ), 
            .I3(n2148), .O(\mult1/n194 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__3202.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__3203 (.I0(\mem_addr[2] ), .I1(\mult1/result[8] ), .I2(\mult_dout[8] ), 
            .I3(n2148), .O(\mult1/n193 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__3203.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__3204 (.I0(\mem_addr[2] ), .I1(\mult1/result[9] ), .I2(\mult_dout[9] ), 
            .I3(n2148), .O(\mult1/n192 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__3204.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__3205 (.I0(\mem_addr[2] ), .I1(\mult1/result[10] ), .I2(\mult_dout[10] ), 
            .I3(n2148), .O(\mult1/n191 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__3205.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__3206 (.I0(\mem_addr[2] ), .I1(\mult1/result[11] ), .I2(\mult_dout[11] ), 
            .I3(n2148), .O(\mult1/n190 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__3206.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__3207 (.I0(\mem_addr[2] ), .I1(\mult1/result[12] ), .I2(\mult_dout[12] ), 
            .I3(n2148), .O(\mult1/n189 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__3207.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__3208 (.I0(\mem_addr[2] ), .I1(\mult1/result[13] ), .I2(\mult_dout[13] ), 
            .I3(n2148), .O(\mult1/n188 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__3208.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__3209 (.I0(\mem_addr[2] ), .I1(\mult1/result[14] ), .I2(\mult_dout[14] ), 
            .I3(n2148), .O(\mult1/n187 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__3209.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__3210 (.I0(\mem_addr[2] ), .I1(\mult1/result[15] ), .I2(\mult_dout[15] ), 
            .I3(n2148), .O(\mult1/n186 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__3210.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__3211 (.I0(\mem_addr[2] ), .I1(\mult1/result[16] ), .I2(\mult_dout[16] ), 
            .I3(n2148), .O(\mult1/n185 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__3211.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__3212 (.I0(\mem_addr[2] ), .I1(\mult1/result[17] ), .I2(\mult_dout[17] ), 
            .I3(n2148), .O(\mult1/n184 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__3212.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__3213 (.I0(\mem_addr[2] ), .I1(\mult1/result[18] ), .I2(\mult_dout[18] ), 
            .I3(n2148), .O(\mult1/n183 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__3213.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__3214 (.I0(\mem_addr[2] ), .I1(\mult1/result[19] ), .I2(\mult_dout[19] ), 
            .I3(n2148), .O(\mult1/n182 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__3214.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__3215 (.I0(\mem_addr[2] ), .I1(\mult1/result[20] ), .I2(\mult_dout[20] ), 
            .I3(n2148), .O(\mult1/n181 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__3215.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__3216 (.I0(\mem_addr[2] ), .I1(\mult1/result[21] ), .I2(\mult_dout[21] ), 
            .I3(n2148), .O(\mult1/n180 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__3216.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__3217 (.I0(\mem_addr[2] ), .I1(\mult1/result[22] ), .I2(\mult_dout[22] ), 
            .I3(n2148), .O(\mult1/n179 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__3217.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__3218 (.I0(\mem_addr[2] ), .I1(\mult1/result[23] ), .I2(\mult_dout[23] ), 
            .I3(n2148), .O(\mult1/n178 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__3218.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__3219 (.I0(\mem_addr[2] ), .I1(\mult1/result[24] ), .I2(\mult_dout[24] ), 
            .I3(n2148), .O(\mult1/n177 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__3219.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__3220 (.I0(\mem_addr[2] ), .I1(\mult1/result[25] ), .I2(\mult_dout[25] ), 
            .I3(n2148), .O(\mult1/n176 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__3220.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__3221 (.I0(\mem_addr[2] ), .I1(\mult1/result[26] ), .I2(\mult_dout[26] ), 
            .I3(n2148), .O(\mult1/n175 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__3221.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__3222 (.I0(\mem_addr[2] ), .I1(\mult1/result[27] ), .I2(\mult_dout[27] ), 
            .I3(n2148), .O(\mult1/n174 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__3222.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__3223 (.I0(\mem_addr[2] ), .I1(\mult1/result[28] ), .I2(\mult_dout[28] ), 
            .I3(n2148), .O(\mult1/n173 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__3223.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__3224 (.I0(\mem_addr[2] ), .I1(\mult1/result[29] ), .I2(\mult_dout[29] ), 
            .I3(n2148), .O(\mult1/n172 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__3224.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__3225 (.I0(\mem_addr[2] ), .I1(\mult1/result[30] ), .I2(\mult_dout[30] ), 
            .I3(n2148), .O(\mult1/n171 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__3225.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__3226 (.I0(\mem_addr[2] ), .I1(\mult1/result[31] ), .I2(\mult_dout[31] ), 
            .I3(n2148), .O(\mult1/n170 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0 */ ;
    defparam LUT__3226.LUTMASK = 16'h44f0;
    EFX_LUT4 LUT__3227 (.I0(\mult1/mult1/state[2] ), .I1(\mult1/mult1/state[1] ), 
            .I2(n209), .O(\mult1/mult1/n132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3227.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3228 (.I0(\mult1/mult1/state[1] ), .I1(\mult1/mult1/state[2] ), 
            .I2(\mult1/mult1/state[0] ), .O(ceg_net913)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9e9e */ ;
    defparam LUT__3228.LUTMASK = 16'h9e9e;
    EFX_LUT4 LUT__3229 (.I0(\mult1/init ), .I1(\mult1/mult1/B[0] ), .I2(\mult1/mult1/state[1] ), 
            .I3(\mult1/mult1/state[0] ), .O(n2149)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__3229.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__3230 (.I0(\mult1/mult1/B[4] ), .I1(\mult1/mult1/B[5] ), 
            .I2(\mult1/mult1/B[6] ), .I3(\mult1/mult1/B[7] ), .O(n2150)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3230.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3231 (.I0(\mult1/mult1/B[1] ), .I1(\mult1/mult1/B[2] ), 
            .I2(\mult1/mult1/B[3] ), .I3(\mult1/mult1/state[1] ), .O(n2151)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__3231.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__3232 (.I0(\mult1/mult1/B[12] ), .I1(\mult1/mult1/B[13] ), 
            .I2(\mult1/mult1/B[14] ), .I3(\mult1/mult1/B[15] ), .O(n2152)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3232.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3233 (.I0(\mult1/mult1/B[8] ), .I1(\mult1/mult1/B[9] ), 
            .I2(\mult1/mult1/B[10] ), .I3(\mult1/mult1/B[11] ), .O(n2153)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3233.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3234 (.I0(n2150), .I1(n2151), .I2(n2152), .I3(n2153), 
            .O(n2154)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3234.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3235 (.I0(n2154), .I1(\mult1/mult1/state[0] ), .I2(\mult1/mult1/state[2] ), 
            .I3(n2149), .O(\mult1/mult1/n64 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__3235.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__3236 (.I0(\mult1/mult1/state[1] ), .I1(\mult1/mult1/state[2] ), 
            .O(ceg_net252)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3236.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3237 (.I0(\mult1/A[0] ), .I1(\mult1/mult1/state[2] ), 
            .O(\mult1/mult1/n81 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3237.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3238 (.I0(\mult1/mult1/state[0] ), .I1(\mult1/mult1/state[2] ), 
            .I2(\mult1/mult1/state[1] ), .O(ceg_net839)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1818 */ ;
    defparam LUT__3238.LUTMASK = 16'h1818;
    EFX_LUT4 LUT__3239 (.I0(\mult1/mult1/B[1] ), .I1(\mult1/B[0] ), .I2(\mult1/mult1/state[2] ), 
            .O(\mult1/mult1/n98 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3239.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3240 (.I0(\mult1/mult1/count[0] ), .I1(\mult1/mult1/state[2] ), 
            .O(\mult1/mult1/n138 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3240.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3241 (.I0(\mult1/mult1/state[0] ), .I1(\mult1/mult1/state[1] ), 
            .I2(resetn), .O(ceg_net847)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__3241.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__3242 (.I0(\mult1/mult1/state[0] ), .I1(\mult1/mult1/state[2] ), 
            .O(\mult1/mult1/n99 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3242.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3243 (.I0(\mult1/mult1/state[0] ), .I1(\mult1/mult1/state[1] ), 
            .I2(\mult1/mult1/state[2] ), .O(ceg_net564)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc2c2 */ ;
    defparam LUT__3243.LUTMASK = 16'hc2c2;
    EFX_LUT4 LUT__3244 (.I0(\mult1/mult1/state[2] ), .I1(\mult1/mult1/state[1] ), 
            .I2(n238), .O(\mult1/mult1/n131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3244.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3245 (.I0(\mult1/mult1/state[2] ), .I1(\mult1/mult1/state[1] ), 
            .I2(n508), .O(\mult1/mult1/n130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3245.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3246 (.I0(\mult1/mult1/state[2] ), .I1(\mult1/mult1/state[1] ), 
            .I2(n506), .O(\mult1/mult1/n129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3246.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3247 (.I0(\mult1/mult1/state[2] ), .I1(\mult1/mult1/state[1] ), 
            .I2(n504), .O(\mult1/mult1/n128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3247.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3248 (.I0(\mult1/mult1/state[2] ), .I1(\mult1/mult1/state[1] ), 
            .I2(n502), .O(\mult1/mult1/n127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3248.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3249 (.I0(\mult1/mult1/state[2] ), .I1(\mult1/mult1/state[1] ), 
            .I2(n500), .O(\mult1/mult1/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3249.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3250 (.I0(\mult1/mult1/state[2] ), .I1(\mult1/mult1/state[1] ), 
            .I2(n498), .O(\mult1/mult1/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3250.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3251 (.I0(\mult1/mult1/state[2] ), .I1(\mult1/mult1/state[1] ), 
            .I2(n496), .O(\mult1/mult1/n124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3251.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3252 (.I0(\mult1/mult1/state[2] ), .I1(\mult1/mult1/state[1] ), 
            .I2(n494), .O(\mult1/mult1/n123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3252.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3253 (.I0(\mult1/mult1/state[2] ), .I1(\mult1/mult1/state[1] ), 
            .I2(n492), .O(\mult1/mult1/n122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3253.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3254 (.I0(\mult1/mult1/state[2] ), .I1(\mult1/mult1/state[1] ), 
            .I2(n490), .O(\mult1/mult1/n121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3254.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3255 (.I0(\mult1/mult1/state[2] ), .I1(\mult1/mult1/state[1] ), 
            .I2(n488), .O(\mult1/mult1/n120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3255.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3256 (.I0(\mult1/mult1/state[2] ), .I1(\mult1/mult1/state[1] ), 
            .I2(n486), .O(\mult1/mult1/n119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3256.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3257 (.I0(\mult1/mult1/state[2] ), .I1(\mult1/mult1/state[1] ), 
            .I2(n484), .O(\mult1/mult1/n118 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3257.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3258 (.I0(\mult1/mult1/state[2] ), .I1(\mult1/mult1/state[1] ), 
            .I2(n482), .O(\mult1/mult1/n117 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3258.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3259 (.I0(\mult1/mult1/state[2] ), .I1(\mult1/mult1/state[1] ), 
            .I2(n480), .O(\mult1/mult1/n116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3259.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3260 (.I0(\mult1/mult1/state[2] ), .I1(\mult1/mult1/state[1] ), 
            .I2(n478), .O(\mult1/mult1/n115 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3260.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3261 (.I0(\mult1/mult1/state[2] ), .I1(\mult1/mult1/state[1] ), 
            .I2(n476), .O(\mult1/mult1/n114 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3261.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3262 (.I0(\mult1/mult1/state[2] ), .I1(\mult1/mult1/state[1] ), 
            .I2(n474), .O(\mult1/mult1/n113 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3262.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3263 (.I0(\mult1/mult1/state[2] ), .I1(\mult1/mult1/state[1] ), 
            .I2(n472), .O(\mult1/mult1/n112 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3263.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3264 (.I0(\mult1/mult1/state[2] ), .I1(\mult1/mult1/state[1] ), 
            .I2(n470), .O(\mult1/mult1/n111 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3264.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3265 (.I0(\mult1/mult1/state[2] ), .I1(\mult1/mult1/state[1] ), 
            .I2(n468), .O(\mult1/mult1/n110 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3265.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3266 (.I0(\mult1/mult1/state[2] ), .I1(\mult1/mult1/state[1] ), 
            .I2(n466), .O(\mult1/mult1/n109 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3266.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3267 (.I0(\mult1/mult1/state[2] ), .I1(\mult1/mult1/state[1] ), 
            .I2(n464), .O(\mult1/mult1/n108 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3267.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3268 (.I0(\mult1/mult1/state[2] ), .I1(\mult1/mult1/state[1] ), 
            .I2(n462), .O(\mult1/mult1/n107 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3268.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3269 (.I0(\mult1/mult1/state[2] ), .I1(\mult1/mult1/state[1] ), 
            .I2(n460), .O(\mult1/mult1/n106 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3269.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3270 (.I0(\mult1/mult1/state[2] ), .I1(\mult1/mult1/state[1] ), 
            .I2(n458), .O(\mult1/mult1/n105 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3270.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3271 (.I0(\mult1/mult1/state[2] ), .I1(\mult1/mult1/state[1] ), 
            .I2(n456), .O(\mult1/mult1/n104 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3271.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3272 (.I0(\mult1/mult1/state[2] ), .I1(\mult1/mult1/state[1] ), 
            .I2(n454), .O(\mult1/mult1/n103 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3272.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3273 (.I0(\mult1/mult1/state[2] ), .I1(\mult1/mult1/state[1] ), 
            .I2(n452), .O(\mult1/mult1/n102 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3273.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3274 (.I0(\mult1/mult1/state[2] ), .I1(\mult1/mult1/state[1] ), 
            .I2(n451), .O(\mult1/mult1/n101 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3274.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3275 (.I0(\mult1/mult1/state[2] ), .I1(\mult1/mult1/state[0] ), 
            .O(\mult1/mult1/n63 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3275.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3276 (.I0(\mult1/mult1/count[0] ), .I1(\mult1/mult1/count[1] ), 
            .I2(\mult1/mult1/state[2] ), .O(\mult1/mult1/n137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__3276.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__3277 (.I0(\mult1/mult1/n137 ), .I1(\mult1/mult1/count[2] ), 
            .I2(\mult1/mult1/count[3] ), .I3(\mult1/mult1/count[4] ), .O(n2155)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3277.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3278 (.I0(\mult1/mult1/state[2] ), .I1(\mult1/init ), 
            .I2(\mult1/mult1/state[1] ), .I3(n2155), .O(n2156)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e */ ;
    defparam LUT__3278.LUTMASK = 16'h000e;
    EFX_LUT4 LUT__3279 (.I0(\mult1/mult1/state[2] ), .I1(n2154), .I2(n2156), 
            .I3(\mult1/mult1/state[0] ), .O(\mult1/mult1/n62 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4 */ ;
    defparam LUT__3279.LUTMASK = 16'h00f4;
    EFX_LUT4 LUT__3280 (.I0(\mult1/mult1/A[0] ), .I1(\mult1/A[1] ), .I2(\mult1/mult1/state[2] ), 
            .O(\mult1/mult1/n80 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3280.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3281 (.I0(\mult1/mult1/A[1] ), .I1(\mult1/A[2] ), .I2(\mult1/mult1/state[2] ), 
            .O(\mult1/mult1/n79 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3281.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3282 (.I0(\mult1/mult1/A[2] ), .I1(\mult1/A[3] ), .I2(\mult1/mult1/state[2] ), 
            .O(\mult1/mult1/n78 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3282.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3283 (.I0(\mult1/mult1/A[3] ), .I1(\mult1/A[4] ), .I2(\mult1/mult1/state[2] ), 
            .O(\mult1/mult1/n77 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3283.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3284 (.I0(\mult1/mult1/A[4] ), .I1(\mult1/A[5] ), .I2(\mult1/mult1/state[2] ), 
            .O(\mult1/mult1/n76 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3284.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3285 (.I0(\mult1/mult1/A[5] ), .I1(\mult1/A[6] ), .I2(\mult1/mult1/state[2] ), 
            .O(\mult1/mult1/n75 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3285.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3286 (.I0(\mult1/mult1/A[6] ), .I1(\mult1/A[7] ), .I2(\mult1/mult1/state[2] ), 
            .O(\mult1/mult1/n74 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3286.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3287 (.I0(\mult1/mult1/A[7] ), .I1(\mult1/A[8] ), .I2(\mult1/mult1/state[2] ), 
            .O(\mult1/mult1/n73 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3287.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3288 (.I0(\mult1/mult1/A[8] ), .I1(\mult1/A[9] ), .I2(\mult1/mult1/state[2] ), 
            .O(\mult1/mult1/n72 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3288.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3289 (.I0(\mult1/mult1/A[9] ), .I1(\mult1/A[10] ), .I2(\mult1/mult1/state[2] ), 
            .O(\mult1/mult1/n71 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3289.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3290 (.I0(\mult1/mult1/A[10] ), .I1(\mult1/A[11] ), .I2(\mult1/mult1/state[2] ), 
            .O(\mult1/mult1/n70 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3290.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3291 (.I0(\mult1/mult1/A[11] ), .I1(\mult1/A[12] ), .I2(\mult1/mult1/state[2] ), 
            .O(\mult1/mult1/n69 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3291.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3292 (.I0(\mult1/mult1/A[12] ), .I1(\mult1/A[13] ), .I2(\mult1/mult1/state[2] ), 
            .O(\mult1/mult1/n68 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3292.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3293 (.I0(\mult1/mult1/A[13] ), .I1(\mult1/A[14] ), .I2(\mult1/mult1/state[2] ), 
            .O(\mult1/mult1/n67 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3293.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3294 (.I0(\mult1/mult1/A[14] ), .I1(\mult1/A[15] ), .I2(\mult1/mult1/state[2] ), 
            .O(\mult1/mult1/n66 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3294.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3295 (.I0(\mult1/mult1/B[2] ), .I1(\mult1/B[1] ), .I2(\mult1/mult1/state[2] ), 
            .O(\mult1/mult1/n97 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3295.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3296 (.I0(\mult1/mult1/B[3] ), .I1(\mult1/B[2] ), .I2(\mult1/mult1/state[2] ), 
            .O(\mult1/mult1/n96 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3296.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3297 (.I0(\mult1/mult1/B[4] ), .I1(\mult1/B[3] ), .I2(\mult1/mult1/state[2] ), 
            .O(\mult1/mult1/n95 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3297.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3298 (.I0(\mult1/mult1/B[5] ), .I1(\mult1/B[4] ), .I2(\mult1/mult1/state[2] ), 
            .O(\mult1/mult1/n94 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3298.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3299 (.I0(\mult1/mult1/B[6] ), .I1(\mult1/B[5] ), .I2(\mult1/mult1/state[2] ), 
            .O(\mult1/mult1/n93 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3299.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3300 (.I0(\mult1/mult1/B[7] ), .I1(\mult1/B[6] ), .I2(\mult1/mult1/state[2] ), 
            .O(\mult1/mult1/n92 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3300.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3301 (.I0(\mult1/mult1/B[8] ), .I1(\mult1/B[7] ), .I2(\mult1/mult1/state[2] ), 
            .O(\mult1/mult1/n91 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3301.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3302 (.I0(\mult1/mult1/B[9] ), .I1(\mult1/B[8] ), .I2(\mult1/mult1/state[2] ), 
            .O(\mult1/mult1/n90 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3302.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3303 (.I0(\mult1/mult1/B[10] ), .I1(\mult1/B[9] ), .I2(\mult1/mult1/state[2] ), 
            .O(\mult1/mult1/n89 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3303.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3304 (.I0(\mult1/mult1/B[11] ), .I1(\mult1/B[10] ), .I2(\mult1/mult1/state[2] ), 
            .O(\mult1/mult1/n88 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3304.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3305 (.I0(\mult1/mult1/B[12] ), .I1(\mult1/B[11] ), .I2(\mult1/mult1/state[2] ), 
            .O(\mult1/mult1/n87 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3305.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3306 (.I0(\mult1/mult1/B[13] ), .I1(\mult1/B[12] ), .I2(\mult1/mult1/state[2] ), 
            .O(\mult1/mult1/n86 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3306.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3307 (.I0(\mult1/mult1/B[14] ), .I1(\mult1/B[13] ), .I2(\mult1/mult1/state[2] ), 
            .O(\mult1/mult1/n85 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3307.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3308 (.I0(\mult1/mult1/B[15] ), .I1(\mult1/B[14] ), .I2(\mult1/mult1/state[2] ), 
            .O(\mult1/mult1/n84 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3308.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3309 (.I0(\mult1/B[15] ), .I1(\mult1/mult1/state[2] ), 
            .O(\mult1/mult1/n83 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3309.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3310 (.I0(\mult1/mult1/count[0] ), .I1(\mult1/mult1/count[1] ), 
            .I2(\mult1/mult1/count[2] ), .I3(\mult1/mult1/state[2] ), .O(\mult1/mult1/n136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;
    defparam LUT__3310.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__3311 (.I0(\mult1/mult1/count[0] ), .I1(\mult1/mult1/count[1] ), 
            .I2(\mult1/mult1/count[2] ), .I3(\mult1/mult1/count[3] ), .O(n2157)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__3311.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__3312 (.I0(n2157), .I1(\mult1/mult1/state[2] ), .O(\mult1/mult1/n135 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3312.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3313 (.I0(\mult1/mult1/count[0] ), .I1(\mult1/mult1/count[1] ), 
            .I2(\mult1/mult1/count[2] ), .I3(\mult1/mult1/count[3] ), .O(n2158)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3313.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3314 (.I0(n2158), .I1(\mult1/mult1/count[4] ), .I2(\mult1/mult1/state[2] ), 
            .O(\mult1/mult1/n134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__3314.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__3315 (.I0(\CPU/instr[24] ), .I1(\CPU/instr[11] ), .I2(\CPU/instr[5] ), 
            .O(n1378)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3315.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3316 (.I0(\CPU/instr[23] ), .I1(\CPU/instr[10] ), .I2(\CPU/instr[5] ), 
            .O(n1381)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3316.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3317 (.I0(\CPU/instr[22] ), .I1(\CPU/instr[9] ), .I2(\CPU/instr[5] ), 
            .O(n1384)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3317.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3318 (.I0(\CPU/instr[21] ), .I1(\CPU/instr[8] ), .I2(\CPU/instr[5] ), 
            .O(n1387)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3318.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3319 (.I0(\CPU/instr[23] ), .I1(\CPU/instr[31] ), .I2(\CPU/instr[3] ), 
            .I3(\CPU/instr[4] ), .O(n1390)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__3319.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__3320 (.I0(\CPU/instr[22] ), .I1(\CPU/instr[31] ), .I2(\CPU/instr[3] ), 
            .I3(\CPU/instr[4] ), .O(n1393)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__3320.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__3321 (.I0(\CPU/instr[21] ), .I1(\CPU/instr[31] ), .I2(\CPU/instr[3] ), 
            .I3(\CPU/instr[4] ), .O(n1396)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__3321.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__3322 (.I0(\CPU/instr[20] ), .I1(\CPU/instr[31] ), .I2(\CPU/instr[3] ), 
            .I3(\CPU/instr[4] ), .O(n1399)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcacc */ ;
    defparam LUT__3322.LUTMASK = 16'hcacc;
    EFX_LUT4 LUT__3323 (.I0(\CPU/instr[31] ), .I1(\CPU/instr[19] ), .I2(\CPU/instr[3] ), 
            .I3(\CPU/instr[4] ), .O(n1402)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca */ ;
    defparam LUT__3323.LUTMASK = 16'hccca;
    EFX_LUT4 LUT__3324 (.I0(\CPU/instr[31] ), .I1(\CPU/instr[18] ), .I2(\CPU/instr[3] ), 
            .I3(\CPU/instr[4] ), .O(n1405)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca */ ;
    defparam LUT__3324.LUTMASK = 16'hccca;
    EFX_LUT4 LUT__3325 (.I0(\CPU/instr[31] ), .I1(\CPU/instr[17] ), .I2(\CPU/instr[3] ), 
            .I3(\CPU/instr[4] ), .O(n1408)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca */ ;
    defparam LUT__3325.LUTMASK = 16'hccca;
    EFX_LUT4 LUT__3326 (.I0(\CPU/instr[31] ), .I1(\CPU/instr[16] ), .I2(\CPU/instr[3] ), 
            .I3(\CPU/instr[4] ), .O(n1411)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca */ ;
    defparam LUT__3326.LUTMASK = 16'hccca;
    EFX_LUT4 LUT__3327 (.I0(\CPU/instr[31] ), .I1(\CPU/instr[15] ), .I2(\CPU/instr[3] ), 
            .I3(\CPU/instr[4] ), .O(n1414)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca */ ;
    defparam LUT__3327.LUTMASK = 16'hccca;
    EFX_LUT4 LUT__3328 (.I0(\CPU/instr[31] ), .I1(\CPU/instr[14] ), .I2(\CPU/instr[3] ), 
            .I3(\CPU/instr[4] ), .O(n1417)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca */ ;
    defparam LUT__3328.LUTMASK = 16'hccca;
    EFX_LUT4 LUT__3329 (.I0(\CPU/instr[31] ), .I1(\CPU/instr[13] ), .I2(\CPU/instr[3] ), 
            .I3(\CPU/instr[4] ), .O(n1420)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca */ ;
    defparam LUT__3329.LUTMASK = 16'hccca;
    EFX_LUT4 LUT__3330 (.I0(\CPU/instr[31] ), .I1(\CPU/instr[12] ), .I2(\CPU/instr[3] ), 
            .I3(\CPU/instr[4] ), .O(n1423)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca */ ;
    defparam LUT__3330.LUTMASK = 16'hccca;
    EFX_LUT4 LUT__3331 (.I0(\CPU/instr[4] ), .I1(\CPU/instr[7] ), .I2(\CPU/instr[20] ), 
            .I3(\CPU/instr[3] ), .O(n1426)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044 */ ;
    defparam LUT__3331.LUTMASK = 16'hf044;
    EFX_LUT4 LUT__3332 (.I0(\CPU/instr[4] ), .I1(\CPU/instr[3] ), .I2(\CPU/instr[30] ), 
            .O(n1429)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__3332.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__3333 (.I0(\CPU/instr[4] ), .I1(\CPU/instr[3] ), .I2(\CPU/instr[29] ), 
            .O(n1432)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__3333.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__3334 (.I0(\CPU/instr[4] ), .I1(\CPU/instr[3] ), .I2(\CPU/instr[28] ), 
            .O(n1435)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__3334.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__3335 (.I0(\CPU/instr[4] ), .I1(\CPU/instr[3] ), .I2(\CPU/instr[27] ), 
            .O(n1438)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__3335.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__3336 (.I0(\CPU/instr[4] ), .I1(\CPU/instr[3] ), .I2(\CPU/instr[26] ), 
            .O(n1441)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__3336.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__3337 (.I0(\CPU/instr[4] ), .I1(\CPU/instr[3] ), .I2(\CPU/instr[25] ), 
            .O(n1444)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__3337.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__3338 (.I0(\CPU/instr[4] ), .I1(\CPU/instr[11] ), .I2(\CPU/instr[24] ), 
            .I3(\CPU/instr[3] ), .O(n1447)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044 */ ;
    defparam LUT__3338.LUTMASK = 16'hf044;
    EFX_LUT4 LUT__3339 (.I0(\CPU/instr[4] ), .I1(\CPU/instr[10] ), .I2(\CPU/instr[23] ), 
            .I3(\CPU/instr[3] ), .O(n1450)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044 */ ;
    defparam LUT__3339.LUTMASK = 16'hf044;
    EFX_LUT4 LUT__3340 (.I0(\CPU/instr[4] ), .I1(\CPU/instr[9] ), .I2(\CPU/instr[22] ), 
            .I3(\CPU/instr[3] ), .O(n1453)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044 */ ;
    defparam LUT__3340.LUTMASK = 16'hf044;
    EFX_LUT4 LUT__2368 (.I0(\mem_rdata[2] ), .I1(\mem_rdata[3] ), .I2(\mem_rdata[5] ), 
            .O(n1589)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__2368.LUTMASK = 16'h1010;
    EFX_GBUFCE CLKBUF__0 (.CE(1'b1), .I(clk), .O(\clk~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__0.CE_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CO__CPU/add_33/i32  (.I0(1'b0), .I1(1'b0), .CI(n2159), 
            .O(n658)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(131)
    defparam \AUX_ADD_CO__CPU/add_33/i32 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CO__CPU/add_33/i32 .I1_POLARITY = 1'b1;
    EFX_FF \CPU/instr[4]~FF_frt_1_frt_2  (.D(n1674), .CE(\CPU/n3447 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/instr[4]~FF_frt_1_frt_2_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/instr[4]~FF_frt_1_frt_2 .CLK_POLARITY = 1'b1;
    defparam \CPU/instr[4]~FF_frt_1_frt_2 .CE_POLARITY = 1'b1;
    defparam \CPU/instr[4]~FF_frt_1_frt_2 .SR_POLARITY = 1'b1;
    defparam \CPU/instr[4]~FF_frt_1_frt_2 .D_POLARITY = 1'b1;
    defparam \CPU/instr[4]~FF_frt_1_frt_2 .SR_SYNC = 1'b1;
    defparam \CPU/instr[4]~FF_frt_1_frt_2 .SR_VALUE = 1'b0;
    defparam \CPU/instr[4]~FF_frt_1_frt_2 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/instr[4]~FF_frt_1  (.D(n1588), .CE(\CPU/n3447 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/instr[4]~FF_frt_1_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/instr[4]~FF_frt_1 .CLK_POLARITY = 1'b1;
    defparam \CPU/instr[4]~FF_frt_1 .CE_POLARITY = 1'b1;
    defparam \CPU/instr[4]~FF_frt_1 .SR_POLARITY = 1'b1;
    defparam \CPU/instr[4]~FF_frt_1 .D_POLARITY = 1'b1;
    defparam \CPU/instr[4]~FF_frt_1 .SR_SYNC = 1'b1;
    defparam \CPU/instr[4]~FF_frt_1 .SR_VALUE = 1'b0;
    defparam \CPU/instr[4]~FF_frt_1 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \CPU/instr[2]~FF_frt_0  (.D(n1589), .CE(\CPU/n3447 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\CPU/instr[2]~FF_frt_0_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // /Work/Proyects/ecb_T8_T113/femtoRV/basic/rtl/cores/cpu/femtorv32_quark.v(369)
    defparam \CPU/instr[2]~FF_frt_0 .CLK_POLARITY = 1'b1;
    defparam \CPU/instr[2]~FF_frt_0 .CE_POLARITY = 1'b1;
    defparam \CPU/instr[2]~FF_frt_0 .SR_POLARITY = 1'b1;
    defparam \CPU/instr[2]~FF_frt_0 .D_POLARITY = 1'b1;
    defparam \CPU/instr[2]~FF_frt_0 .SR_SYNC = 1'b1;
    defparam \CPU/instr[2]~FF_frt_0 .SR_VALUE = 1'b0;
    defparam \CPU/instr[2]~FF_frt_0 .SR_SYNC_PRIORITY = 1'b1;
    
endmodule

//
// Verific Verilog Description of module EFX_FF_2b382480_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_2b382480_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_2b382480_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_2b382480_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_2b382480_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_2b382480_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_2b382480_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_2b382480_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_2b382480_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_2b382480_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_2b382480_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_2b382480_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b382480__1_1_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b382480__16_16_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b382480__16_16_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b382480__16_16_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b382480__16_16_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b382480__1_1_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b382480__1_1_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b382480__1_1_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b382480__1_1_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b382480__1_1_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b382480__1_1_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b382480__1_1_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b382480__1_1_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b382480__1_1_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b382480__1_1_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b382480__1_1_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b382480__1_1_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b382480__1_1_17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b382480__1_1_18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b382480__1_1_19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b382480__1_1_20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b382480__1_1_21
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b382480__1_1_22
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b382480__1_1_23
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b382480__1_1_24
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b382480__1_1_25
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b382480__1_1_26
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b382480__1_1_27
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b382480__1_1_28
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b382480__1_1_29
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b382480__1_1_30
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b382480__1_1_31
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b382480__1_1_32
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b382480__1_1_33
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b382480__1_1_34
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_2b382480__1_1_35
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_21
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_22
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_23
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_24
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_25
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_26
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_27
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_28
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_29
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_30
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_31
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_32
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_33
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_34
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_35
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_36
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_37
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_38
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_39
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_40
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_41
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_42
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_43
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_44
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_45
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_46
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_47
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_48
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_49
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_50
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_51
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_52
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_53
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_54
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_55
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_56
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_57
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_58
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_59
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_60
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_61
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_62
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_63
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_64
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_65
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_66
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_67
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_68
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_69
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_70
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_71
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_72
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_73
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_74
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_75
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_76
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_77
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_78
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_79
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_80
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_81
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_82
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_83
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_84
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_85
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_86
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_87
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_88
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_89
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_90
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_91
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_92
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_93
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_94
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_95
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_96
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_97
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_98
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_99
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_100
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_101
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_102
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_103
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_104
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_105
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_106
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_107
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_108
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_109
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_110
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_111
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_112
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_113
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_114
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_115
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_116
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_117
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_118
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_119
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_120
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_121
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_122
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_123
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_124
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_125
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_126
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_127
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_128
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_129
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_130
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_131
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_2b382480_132
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_GBUFCE_2b382480_0
// module not written out since it is a black box. 
//

